library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- library SYSTEM_TYPES;
use work.SYSTEM_TYPES.ALL;

-- library CUSTOM_TYPES;
use work.CUSTOM_TYPES.ALL;

-- User defined packages here
-- #### USER-DATA-IMPORTS-START
-- #### USER-DATA-IMPORTS-END

entity Decoder_n_Bit is
  port(


    -- Top-level bus DecoderInput_0 signals
    DecoderInput_0_Value: in T_SYSTEM_BOOL;

    -- Top-level bus DecoderNOTInput_0 signals
    DecoderNOTInput_0_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderInput_1 signals
    DecoderInput_1_Value: in T_SYSTEM_BOOL;

    -- Top-level bus DecoderNOTInput_1 signals
    DecoderNOTInput_1_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderInput_2 signals
    DecoderInput_2_Value: in T_SYSTEM_BOOL;

    -- Top-level bus DecoderNOTInput_2 signals
    DecoderNOTInput_2_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderInput_3 signals
    DecoderInput_3_Value: in T_SYSTEM_BOOL;

    -- Top-level bus DecoderNOTInput_3 signals
    DecoderNOTInput_3_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderInput_4 signals
    DecoderInput_4_Value: in T_SYSTEM_BOOL;

    -- Top-level bus DecoderNOTInput_4 signals
    DecoderNOTInput_4_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderInput_5 signals
    DecoderInput_5_Value: in T_SYSTEM_BOOL;

    -- Top-level bus DecoderNOTInput_5 signals
    DecoderNOTInput_5_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderInput_6 signals
    DecoderInput_6_Value: in T_SYSTEM_BOOL;

    -- Top-level bus DecoderNOTInput_6 signals
    DecoderNOTInput_6_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderInput_7 signals
    DecoderInput_7_Value: in T_SYSTEM_BOOL;

    -- Top-level bus DecoderNOTInput_7 signals
    DecoderNOTInput_7_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_0 signals
    DecoderOutput_0_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_1 signals
    DecoderOutput_1_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_2 signals
    DecoderOutput_2_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_3 signals
    DecoderOutput_3_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_4 signals
    DecoderOutput_4_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_5 signals
    DecoderOutput_5_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_6 signals
    DecoderOutput_6_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_7 signals
    DecoderOutput_7_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_8 signals
    DecoderOutput_8_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_9 signals
    DecoderOutput_9_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_10 signals
    DecoderOutput_10_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_11 signals
    DecoderOutput_11_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_12 signals
    DecoderOutput_12_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_13 signals
    DecoderOutput_13_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_14 signals
    DecoderOutput_14_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_15 signals
    DecoderOutput_15_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_16 signals
    DecoderOutput_16_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_17 signals
    DecoderOutput_17_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_18 signals
    DecoderOutput_18_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_19 signals
    DecoderOutput_19_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_20 signals
    DecoderOutput_20_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_21 signals
    DecoderOutput_21_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_22 signals
    DecoderOutput_22_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_23 signals
    DecoderOutput_23_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_24 signals
    DecoderOutput_24_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_25 signals
    DecoderOutput_25_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_26 signals
    DecoderOutput_26_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_27 signals
    DecoderOutput_27_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_28 signals
    DecoderOutput_28_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_29 signals
    DecoderOutput_29_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_30 signals
    DecoderOutput_30_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_31 signals
    DecoderOutput_31_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_32 signals
    DecoderOutput_32_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_33 signals
    DecoderOutput_33_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_34 signals
    DecoderOutput_34_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_35 signals
    DecoderOutput_35_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_36 signals
    DecoderOutput_36_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_37 signals
    DecoderOutput_37_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_38 signals
    DecoderOutput_38_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_39 signals
    DecoderOutput_39_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_40 signals
    DecoderOutput_40_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_41 signals
    DecoderOutput_41_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_42 signals
    DecoderOutput_42_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_43 signals
    DecoderOutput_43_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_44 signals
    DecoderOutput_44_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_45 signals
    DecoderOutput_45_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_46 signals
    DecoderOutput_46_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_47 signals
    DecoderOutput_47_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_48 signals
    DecoderOutput_48_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_49 signals
    DecoderOutput_49_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_50 signals
    DecoderOutput_50_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_51 signals
    DecoderOutput_51_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_52 signals
    DecoderOutput_52_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_53 signals
    DecoderOutput_53_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_54 signals
    DecoderOutput_54_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_55 signals
    DecoderOutput_55_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_56 signals
    DecoderOutput_56_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_57 signals
    DecoderOutput_57_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_58 signals
    DecoderOutput_58_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_59 signals
    DecoderOutput_59_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_60 signals
    DecoderOutput_60_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_61 signals
    DecoderOutput_61_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_62 signals
    DecoderOutput_62_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_63 signals
    DecoderOutput_63_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_64 signals
    DecoderOutput_64_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_65 signals
    DecoderOutput_65_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_66 signals
    DecoderOutput_66_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_67 signals
    DecoderOutput_67_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_68 signals
    DecoderOutput_68_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_69 signals
    DecoderOutput_69_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_70 signals
    DecoderOutput_70_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_71 signals
    DecoderOutput_71_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_72 signals
    DecoderOutput_72_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_73 signals
    DecoderOutput_73_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_74 signals
    DecoderOutput_74_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_75 signals
    DecoderOutput_75_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_76 signals
    DecoderOutput_76_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_77 signals
    DecoderOutput_77_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_78 signals
    DecoderOutput_78_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_79 signals
    DecoderOutput_79_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_80 signals
    DecoderOutput_80_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_81 signals
    DecoderOutput_81_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_82 signals
    DecoderOutput_82_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_83 signals
    DecoderOutput_83_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_84 signals
    DecoderOutput_84_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_85 signals
    DecoderOutput_85_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_86 signals
    DecoderOutput_86_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_87 signals
    DecoderOutput_87_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_88 signals
    DecoderOutput_88_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_89 signals
    DecoderOutput_89_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_90 signals
    DecoderOutput_90_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_91 signals
    DecoderOutput_91_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_92 signals
    DecoderOutput_92_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_93 signals
    DecoderOutput_93_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_94 signals
    DecoderOutput_94_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_95 signals
    DecoderOutput_95_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_96 signals
    DecoderOutput_96_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_97 signals
    DecoderOutput_97_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_98 signals
    DecoderOutput_98_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_99 signals
    DecoderOutput_99_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_100 signals
    DecoderOutput_100_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_101 signals
    DecoderOutput_101_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_102 signals
    DecoderOutput_102_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_103 signals
    DecoderOutput_103_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_104 signals
    DecoderOutput_104_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_105 signals
    DecoderOutput_105_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_106 signals
    DecoderOutput_106_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_107 signals
    DecoderOutput_107_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_108 signals
    DecoderOutput_108_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_109 signals
    DecoderOutput_109_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_110 signals
    DecoderOutput_110_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_111 signals
    DecoderOutput_111_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_112 signals
    DecoderOutput_112_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_113 signals
    DecoderOutput_113_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_114 signals
    DecoderOutput_114_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_115 signals
    DecoderOutput_115_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_116 signals
    DecoderOutput_116_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_117 signals
    DecoderOutput_117_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_118 signals
    DecoderOutput_118_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_119 signals
    DecoderOutput_119_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_120 signals
    DecoderOutput_120_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_121 signals
    DecoderOutput_121_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_122 signals
    DecoderOutput_122_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_123 signals
    DecoderOutput_123_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_124 signals
    DecoderOutput_124_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_125 signals
    DecoderOutput_125_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_126 signals
    DecoderOutput_126_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_127 signals
    DecoderOutput_127_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_128 signals
    DecoderOutput_128_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_129 signals
    DecoderOutput_129_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_130 signals
    DecoderOutput_130_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_131 signals
    DecoderOutput_131_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_132 signals
    DecoderOutput_132_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_133 signals
    DecoderOutput_133_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_134 signals
    DecoderOutput_134_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_135 signals
    DecoderOutput_135_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_136 signals
    DecoderOutput_136_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_137 signals
    DecoderOutput_137_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_138 signals
    DecoderOutput_138_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_139 signals
    DecoderOutput_139_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_140 signals
    DecoderOutput_140_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_141 signals
    DecoderOutput_141_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_142 signals
    DecoderOutput_142_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_143 signals
    DecoderOutput_143_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_144 signals
    DecoderOutput_144_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_145 signals
    DecoderOutput_145_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_146 signals
    DecoderOutput_146_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_147 signals
    DecoderOutput_147_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_148 signals
    DecoderOutput_148_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_149 signals
    DecoderOutput_149_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_150 signals
    DecoderOutput_150_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_151 signals
    DecoderOutput_151_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_152 signals
    DecoderOutput_152_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_153 signals
    DecoderOutput_153_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_154 signals
    DecoderOutput_154_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_155 signals
    DecoderOutput_155_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_156 signals
    DecoderOutput_156_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_157 signals
    DecoderOutput_157_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_158 signals
    DecoderOutput_158_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_159 signals
    DecoderOutput_159_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_160 signals
    DecoderOutput_160_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_161 signals
    DecoderOutput_161_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_162 signals
    DecoderOutput_162_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_163 signals
    DecoderOutput_163_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_164 signals
    DecoderOutput_164_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_165 signals
    DecoderOutput_165_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_166 signals
    DecoderOutput_166_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_167 signals
    DecoderOutput_167_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_168 signals
    DecoderOutput_168_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_169 signals
    DecoderOutput_169_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_170 signals
    DecoderOutput_170_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_171 signals
    DecoderOutput_171_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_172 signals
    DecoderOutput_172_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_173 signals
    DecoderOutput_173_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_174 signals
    DecoderOutput_174_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_175 signals
    DecoderOutput_175_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_176 signals
    DecoderOutput_176_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_177 signals
    DecoderOutput_177_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_178 signals
    DecoderOutput_178_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_179 signals
    DecoderOutput_179_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_180 signals
    DecoderOutput_180_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_181 signals
    DecoderOutput_181_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_182 signals
    DecoderOutput_182_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_183 signals
    DecoderOutput_183_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_184 signals
    DecoderOutput_184_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_185 signals
    DecoderOutput_185_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_186 signals
    DecoderOutput_186_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_187 signals
    DecoderOutput_187_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_188 signals
    DecoderOutput_188_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_189 signals
    DecoderOutput_189_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_190 signals
    DecoderOutput_190_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_191 signals
    DecoderOutput_191_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_192 signals
    DecoderOutput_192_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_193 signals
    DecoderOutput_193_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_194 signals
    DecoderOutput_194_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_195 signals
    DecoderOutput_195_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_196 signals
    DecoderOutput_196_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_197 signals
    DecoderOutput_197_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_198 signals
    DecoderOutput_198_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_199 signals
    DecoderOutput_199_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_200 signals
    DecoderOutput_200_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_201 signals
    DecoderOutput_201_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_202 signals
    DecoderOutput_202_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_203 signals
    DecoderOutput_203_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_204 signals
    DecoderOutput_204_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_205 signals
    DecoderOutput_205_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_206 signals
    DecoderOutput_206_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_207 signals
    DecoderOutput_207_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_208 signals
    DecoderOutput_208_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_209 signals
    DecoderOutput_209_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_210 signals
    DecoderOutput_210_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_211 signals
    DecoderOutput_211_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_212 signals
    DecoderOutput_212_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_213 signals
    DecoderOutput_213_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_214 signals
    DecoderOutput_214_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_215 signals
    DecoderOutput_215_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_216 signals
    DecoderOutput_216_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_217 signals
    DecoderOutput_217_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_218 signals
    DecoderOutput_218_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_219 signals
    DecoderOutput_219_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_220 signals
    DecoderOutput_220_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_221 signals
    DecoderOutput_221_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_222 signals
    DecoderOutput_222_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_223 signals
    DecoderOutput_223_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_224 signals
    DecoderOutput_224_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_225 signals
    DecoderOutput_225_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_226 signals
    DecoderOutput_226_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_227 signals
    DecoderOutput_227_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_228 signals
    DecoderOutput_228_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_229 signals
    DecoderOutput_229_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_230 signals
    DecoderOutput_230_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_231 signals
    DecoderOutput_231_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_232 signals
    DecoderOutput_232_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_233 signals
    DecoderOutput_233_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_234 signals
    DecoderOutput_234_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_235 signals
    DecoderOutput_235_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_236 signals
    DecoderOutput_236_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_237 signals
    DecoderOutput_237_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_238 signals
    DecoderOutput_238_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_239 signals
    DecoderOutput_239_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_240 signals
    DecoderOutput_240_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_241 signals
    DecoderOutput_241_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_242 signals
    DecoderOutput_242_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_243 signals
    DecoderOutput_243_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_244 signals
    DecoderOutput_244_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_245 signals
    DecoderOutput_245_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_246 signals
    DecoderOutput_246_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_247 signals
    DecoderOutput_247_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_248 signals
    DecoderOutput_248_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_249 signals
    DecoderOutput_249_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_250 signals
    DecoderOutput_250_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_251 signals
    DecoderOutput_251_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_252 signals
    DecoderOutput_252_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_253 signals
    DecoderOutput_253_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_254 signals
    DecoderOutput_254_Value: out T_SYSTEM_BOOL;

    -- Top-level bus DecoderOutput_255 signals
    DecoderOutput_255_Value: out T_SYSTEM_BOOL;



    -- User defined signals here
    -- #### USER-DATA-ENTITYSIGNALS-START
    -- #### USER-DATA-ENTITYSIGNALS-END

    -- Enable signal
    ENB : in Std_logic;

    -- Finished signal
    FIN : out Std_logic;

	-- Reset signal
    RST : in Std_logic;

	-- Clock signal
	CLK : in Std_logic
  );
end Decoder_n_Bit;

architecture RTL of Decoder_n_Bit is  
    -- User defined signals here
    -- #### USER-DATA-SIGNALS-START
    -- #### USER-DATA-SIGNALS-END


    -- Process ready triggers

    signal FIN_NOTGate_0, RDY_NOTGate_0 : std_logic;

    signal FIN_NOTGate_1, RDY_NOTGate_1 : std_logic;

    signal FIN_NOTGate_2, RDY_NOTGate_2 : std_logic;

    signal FIN_NOTGate_3, RDY_NOTGate_3 : std_logic;

    signal FIN_NOTGate_4, RDY_NOTGate_4 : std_logic;

    signal FIN_NOTGate_5, RDY_NOTGate_5 : std_logic;

    signal FIN_NOTGate_6, RDY_NOTGate_6 : std_logic;

    signal FIN_NOTGate_7, RDY_NOTGate_7 : std_logic;

    signal FIN_ANDGate_0, RDY_ANDGate_0 : std_logic;

    signal FIN_ANDGate_1, RDY_ANDGate_1 : std_logic;

    signal FIN_ANDGate_2, RDY_ANDGate_2 : std_logic;

    signal FIN_ANDGate_3, RDY_ANDGate_3 : std_logic;

    signal FIN_ANDGate_4, RDY_ANDGate_4 : std_logic;

    signal FIN_ANDGate_5, RDY_ANDGate_5 : std_logic;

    signal FIN_ANDGate_6, RDY_ANDGate_6 : std_logic;

    signal FIN_ANDGate_7, RDY_ANDGate_7 : std_logic;

    signal FIN_ANDGate_8, RDY_ANDGate_8 : std_logic;

    signal FIN_ANDGate_9, RDY_ANDGate_9 : std_logic;

    signal FIN_ANDGate_10, RDY_ANDGate_10 : std_logic;

    signal FIN_ANDGate_11, RDY_ANDGate_11 : std_logic;

    signal FIN_ANDGate_12, RDY_ANDGate_12 : std_logic;

    signal FIN_ANDGate_13, RDY_ANDGate_13 : std_logic;

    signal FIN_ANDGate_14, RDY_ANDGate_14 : std_logic;

    signal FIN_ANDGate_15, RDY_ANDGate_15 : std_logic;

    signal FIN_ANDGate_16, RDY_ANDGate_16 : std_logic;

    signal FIN_ANDGate_17, RDY_ANDGate_17 : std_logic;

    signal FIN_ANDGate_18, RDY_ANDGate_18 : std_logic;

    signal FIN_ANDGate_19, RDY_ANDGate_19 : std_logic;

    signal FIN_ANDGate_20, RDY_ANDGate_20 : std_logic;

    signal FIN_ANDGate_21, RDY_ANDGate_21 : std_logic;

    signal FIN_ANDGate_22, RDY_ANDGate_22 : std_logic;

    signal FIN_ANDGate_23, RDY_ANDGate_23 : std_logic;

    signal FIN_ANDGate_24, RDY_ANDGate_24 : std_logic;

    signal FIN_ANDGate_25, RDY_ANDGate_25 : std_logic;

    signal FIN_ANDGate_26, RDY_ANDGate_26 : std_logic;

    signal FIN_ANDGate_27, RDY_ANDGate_27 : std_logic;

    signal FIN_ANDGate_28, RDY_ANDGate_28 : std_logic;

    signal FIN_ANDGate_29, RDY_ANDGate_29 : std_logic;

    signal FIN_ANDGate_30, RDY_ANDGate_30 : std_logic;

    signal FIN_ANDGate_31, RDY_ANDGate_31 : std_logic;

    signal FIN_ANDGate_32, RDY_ANDGate_32 : std_logic;

    signal FIN_ANDGate_33, RDY_ANDGate_33 : std_logic;

    signal FIN_ANDGate_34, RDY_ANDGate_34 : std_logic;

    signal FIN_ANDGate_35, RDY_ANDGate_35 : std_logic;

    signal FIN_ANDGate_36, RDY_ANDGate_36 : std_logic;

    signal FIN_ANDGate_37, RDY_ANDGate_37 : std_logic;

    signal FIN_ANDGate_38, RDY_ANDGate_38 : std_logic;

    signal FIN_ANDGate_39, RDY_ANDGate_39 : std_logic;

    signal FIN_ANDGate_40, RDY_ANDGate_40 : std_logic;

    signal FIN_ANDGate_41, RDY_ANDGate_41 : std_logic;

    signal FIN_ANDGate_42, RDY_ANDGate_42 : std_logic;

    signal FIN_ANDGate_43, RDY_ANDGate_43 : std_logic;

    signal FIN_ANDGate_44, RDY_ANDGate_44 : std_logic;

    signal FIN_ANDGate_45, RDY_ANDGate_45 : std_logic;

    signal FIN_ANDGate_46, RDY_ANDGate_46 : std_logic;

    signal FIN_ANDGate_47, RDY_ANDGate_47 : std_logic;

    signal FIN_ANDGate_48, RDY_ANDGate_48 : std_logic;

    signal FIN_ANDGate_49, RDY_ANDGate_49 : std_logic;

    signal FIN_ANDGate_50, RDY_ANDGate_50 : std_logic;

    signal FIN_ANDGate_51, RDY_ANDGate_51 : std_logic;

    signal FIN_ANDGate_52, RDY_ANDGate_52 : std_logic;

    signal FIN_ANDGate_53, RDY_ANDGate_53 : std_logic;

    signal FIN_ANDGate_54, RDY_ANDGate_54 : std_logic;

    signal FIN_ANDGate_55, RDY_ANDGate_55 : std_logic;

    signal FIN_ANDGate_56, RDY_ANDGate_56 : std_logic;

    signal FIN_ANDGate_57, RDY_ANDGate_57 : std_logic;

    signal FIN_ANDGate_58, RDY_ANDGate_58 : std_logic;

    signal FIN_ANDGate_59, RDY_ANDGate_59 : std_logic;

    signal FIN_ANDGate_60, RDY_ANDGate_60 : std_logic;

    signal FIN_ANDGate_61, RDY_ANDGate_61 : std_logic;

    signal FIN_ANDGate_62, RDY_ANDGate_62 : std_logic;

    signal FIN_ANDGate_63, RDY_ANDGate_63 : std_logic;

    signal FIN_ANDGate_64, RDY_ANDGate_64 : std_logic;

    signal FIN_ANDGate_65, RDY_ANDGate_65 : std_logic;

    signal FIN_ANDGate_66, RDY_ANDGate_66 : std_logic;

    signal FIN_ANDGate_67, RDY_ANDGate_67 : std_logic;

    signal FIN_ANDGate_68, RDY_ANDGate_68 : std_logic;

    signal FIN_ANDGate_69, RDY_ANDGate_69 : std_logic;

    signal FIN_ANDGate_70, RDY_ANDGate_70 : std_logic;

    signal FIN_ANDGate_71, RDY_ANDGate_71 : std_logic;

    signal FIN_ANDGate_72, RDY_ANDGate_72 : std_logic;

    signal FIN_ANDGate_73, RDY_ANDGate_73 : std_logic;

    signal FIN_ANDGate_74, RDY_ANDGate_74 : std_logic;

    signal FIN_ANDGate_75, RDY_ANDGate_75 : std_logic;

    signal FIN_ANDGate_76, RDY_ANDGate_76 : std_logic;

    signal FIN_ANDGate_77, RDY_ANDGate_77 : std_logic;

    signal FIN_ANDGate_78, RDY_ANDGate_78 : std_logic;

    signal FIN_ANDGate_79, RDY_ANDGate_79 : std_logic;

    signal FIN_ANDGate_80, RDY_ANDGate_80 : std_logic;

    signal FIN_ANDGate_81, RDY_ANDGate_81 : std_logic;

    signal FIN_ANDGate_82, RDY_ANDGate_82 : std_logic;

    signal FIN_ANDGate_83, RDY_ANDGate_83 : std_logic;

    signal FIN_ANDGate_84, RDY_ANDGate_84 : std_logic;

    signal FIN_ANDGate_85, RDY_ANDGate_85 : std_logic;

    signal FIN_ANDGate_86, RDY_ANDGate_86 : std_logic;

    signal FIN_ANDGate_87, RDY_ANDGate_87 : std_logic;

    signal FIN_ANDGate_88, RDY_ANDGate_88 : std_logic;

    signal FIN_ANDGate_89, RDY_ANDGate_89 : std_logic;

    signal FIN_ANDGate_90, RDY_ANDGate_90 : std_logic;

    signal FIN_ANDGate_91, RDY_ANDGate_91 : std_logic;

    signal FIN_ANDGate_92, RDY_ANDGate_92 : std_logic;

    signal FIN_ANDGate_93, RDY_ANDGate_93 : std_logic;

    signal FIN_ANDGate_94, RDY_ANDGate_94 : std_logic;

    signal FIN_ANDGate_95, RDY_ANDGate_95 : std_logic;

    signal FIN_ANDGate_96, RDY_ANDGate_96 : std_logic;

    signal FIN_ANDGate_97, RDY_ANDGate_97 : std_logic;

    signal FIN_ANDGate_98, RDY_ANDGate_98 : std_logic;

    signal FIN_ANDGate_99, RDY_ANDGate_99 : std_logic;

    signal FIN_ANDGate_100, RDY_ANDGate_100 : std_logic;

    signal FIN_ANDGate_101, RDY_ANDGate_101 : std_logic;

    signal FIN_ANDGate_102, RDY_ANDGate_102 : std_logic;

    signal FIN_ANDGate_103, RDY_ANDGate_103 : std_logic;

    signal FIN_ANDGate_104, RDY_ANDGate_104 : std_logic;

    signal FIN_ANDGate_105, RDY_ANDGate_105 : std_logic;

    signal FIN_ANDGate_106, RDY_ANDGate_106 : std_logic;

    signal FIN_ANDGate_107, RDY_ANDGate_107 : std_logic;

    signal FIN_ANDGate_108, RDY_ANDGate_108 : std_logic;

    signal FIN_ANDGate_109, RDY_ANDGate_109 : std_logic;

    signal FIN_ANDGate_110, RDY_ANDGate_110 : std_logic;

    signal FIN_ANDGate_111, RDY_ANDGate_111 : std_logic;

    signal FIN_ANDGate_112, RDY_ANDGate_112 : std_logic;

    signal FIN_ANDGate_113, RDY_ANDGate_113 : std_logic;

    signal FIN_ANDGate_114, RDY_ANDGate_114 : std_logic;

    signal FIN_ANDGate_115, RDY_ANDGate_115 : std_logic;

    signal FIN_ANDGate_116, RDY_ANDGate_116 : std_logic;

    signal FIN_ANDGate_117, RDY_ANDGate_117 : std_logic;

    signal FIN_ANDGate_118, RDY_ANDGate_118 : std_logic;

    signal FIN_ANDGate_119, RDY_ANDGate_119 : std_logic;

    signal FIN_ANDGate_120, RDY_ANDGate_120 : std_logic;

    signal FIN_ANDGate_121, RDY_ANDGate_121 : std_logic;

    signal FIN_ANDGate_122, RDY_ANDGate_122 : std_logic;

    signal FIN_ANDGate_123, RDY_ANDGate_123 : std_logic;

    signal FIN_ANDGate_124, RDY_ANDGate_124 : std_logic;

    signal FIN_ANDGate_125, RDY_ANDGate_125 : std_logic;

    signal FIN_ANDGate_126, RDY_ANDGate_126 : std_logic;

    signal FIN_ANDGate_127, RDY_ANDGate_127 : std_logic;

    signal FIN_ANDGate_128, RDY_ANDGate_128 : std_logic;

    signal FIN_ANDGate_129, RDY_ANDGate_129 : std_logic;

    signal FIN_ANDGate_130, RDY_ANDGate_130 : std_logic;

    signal FIN_ANDGate_131, RDY_ANDGate_131 : std_logic;

    signal FIN_ANDGate_132, RDY_ANDGate_132 : std_logic;

    signal FIN_ANDGate_133, RDY_ANDGate_133 : std_logic;

    signal FIN_ANDGate_134, RDY_ANDGate_134 : std_logic;

    signal FIN_ANDGate_135, RDY_ANDGate_135 : std_logic;

    signal FIN_ANDGate_136, RDY_ANDGate_136 : std_logic;

    signal FIN_ANDGate_137, RDY_ANDGate_137 : std_logic;

    signal FIN_ANDGate_138, RDY_ANDGate_138 : std_logic;

    signal FIN_ANDGate_139, RDY_ANDGate_139 : std_logic;

    signal FIN_ANDGate_140, RDY_ANDGate_140 : std_logic;

    signal FIN_ANDGate_141, RDY_ANDGate_141 : std_logic;

    signal FIN_ANDGate_142, RDY_ANDGate_142 : std_logic;

    signal FIN_ANDGate_143, RDY_ANDGate_143 : std_logic;

    signal FIN_ANDGate_144, RDY_ANDGate_144 : std_logic;

    signal FIN_ANDGate_145, RDY_ANDGate_145 : std_logic;

    signal FIN_ANDGate_146, RDY_ANDGate_146 : std_logic;

    signal FIN_ANDGate_147, RDY_ANDGate_147 : std_logic;

    signal FIN_ANDGate_148, RDY_ANDGate_148 : std_logic;

    signal FIN_ANDGate_149, RDY_ANDGate_149 : std_logic;

    signal FIN_ANDGate_150, RDY_ANDGate_150 : std_logic;

    signal FIN_ANDGate_151, RDY_ANDGate_151 : std_logic;

    signal FIN_ANDGate_152, RDY_ANDGate_152 : std_logic;

    signal FIN_ANDGate_153, RDY_ANDGate_153 : std_logic;

    signal FIN_ANDGate_154, RDY_ANDGate_154 : std_logic;

    signal FIN_ANDGate_155, RDY_ANDGate_155 : std_logic;

    signal FIN_ANDGate_156, RDY_ANDGate_156 : std_logic;

    signal FIN_ANDGate_157, RDY_ANDGate_157 : std_logic;

    signal FIN_ANDGate_158, RDY_ANDGate_158 : std_logic;

    signal FIN_ANDGate_159, RDY_ANDGate_159 : std_logic;

    signal FIN_ANDGate_160, RDY_ANDGate_160 : std_logic;

    signal FIN_ANDGate_161, RDY_ANDGate_161 : std_logic;

    signal FIN_ANDGate_162, RDY_ANDGate_162 : std_logic;

    signal FIN_ANDGate_163, RDY_ANDGate_163 : std_logic;

    signal FIN_ANDGate_164, RDY_ANDGate_164 : std_logic;

    signal FIN_ANDGate_165, RDY_ANDGate_165 : std_logic;

    signal FIN_ANDGate_166, RDY_ANDGate_166 : std_logic;

    signal FIN_ANDGate_167, RDY_ANDGate_167 : std_logic;

    signal FIN_ANDGate_168, RDY_ANDGate_168 : std_logic;

    signal FIN_ANDGate_169, RDY_ANDGate_169 : std_logic;

    signal FIN_ANDGate_170, RDY_ANDGate_170 : std_logic;

    signal FIN_ANDGate_171, RDY_ANDGate_171 : std_logic;

    signal FIN_ANDGate_172, RDY_ANDGate_172 : std_logic;

    signal FIN_ANDGate_173, RDY_ANDGate_173 : std_logic;

    signal FIN_ANDGate_174, RDY_ANDGate_174 : std_logic;

    signal FIN_ANDGate_175, RDY_ANDGate_175 : std_logic;

    signal FIN_ANDGate_176, RDY_ANDGate_176 : std_logic;

    signal FIN_ANDGate_177, RDY_ANDGate_177 : std_logic;

    signal FIN_ANDGate_178, RDY_ANDGate_178 : std_logic;

    signal FIN_ANDGate_179, RDY_ANDGate_179 : std_logic;

    signal FIN_ANDGate_180, RDY_ANDGate_180 : std_logic;

    signal FIN_ANDGate_181, RDY_ANDGate_181 : std_logic;

    signal FIN_ANDGate_182, RDY_ANDGate_182 : std_logic;

    signal FIN_ANDGate_183, RDY_ANDGate_183 : std_logic;

    signal FIN_ANDGate_184, RDY_ANDGate_184 : std_logic;

    signal FIN_ANDGate_185, RDY_ANDGate_185 : std_logic;

    signal FIN_ANDGate_186, RDY_ANDGate_186 : std_logic;

    signal FIN_ANDGate_187, RDY_ANDGate_187 : std_logic;

    signal FIN_ANDGate_188, RDY_ANDGate_188 : std_logic;

    signal FIN_ANDGate_189, RDY_ANDGate_189 : std_logic;

    signal FIN_ANDGate_190, RDY_ANDGate_190 : std_logic;

    signal FIN_ANDGate_191, RDY_ANDGate_191 : std_logic;

    signal FIN_ANDGate_192, RDY_ANDGate_192 : std_logic;

    signal FIN_ANDGate_193, RDY_ANDGate_193 : std_logic;

    signal FIN_ANDGate_194, RDY_ANDGate_194 : std_logic;

    signal FIN_ANDGate_195, RDY_ANDGate_195 : std_logic;

    signal FIN_ANDGate_196, RDY_ANDGate_196 : std_logic;

    signal FIN_ANDGate_197, RDY_ANDGate_197 : std_logic;

    signal FIN_ANDGate_198, RDY_ANDGate_198 : std_logic;

    signal FIN_ANDGate_199, RDY_ANDGate_199 : std_logic;

    signal FIN_ANDGate_200, RDY_ANDGate_200 : std_logic;

    signal FIN_ANDGate_201, RDY_ANDGate_201 : std_logic;

    signal FIN_ANDGate_202, RDY_ANDGate_202 : std_logic;

    signal FIN_ANDGate_203, RDY_ANDGate_203 : std_logic;

    signal FIN_ANDGate_204, RDY_ANDGate_204 : std_logic;

    signal FIN_ANDGate_205, RDY_ANDGate_205 : std_logic;

    signal FIN_ANDGate_206, RDY_ANDGate_206 : std_logic;

    signal FIN_ANDGate_207, RDY_ANDGate_207 : std_logic;

    signal FIN_ANDGate_208, RDY_ANDGate_208 : std_logic;

    signal FIN_ANDGate_209, RDY_ANDGate_209 : std_logic;

    signal FIN_ANDGate_210, RDY_ANDGate_210 : std_logic;

    signal FIN_ANDGate_211, RDY_ANDGate_211 : std_logic;

    signal FIN_ANDGate_212, RDY_ANDGate_212 : std_logic;

    signal FIN_ANDGate_213, RDY_ANDGate_213 : std_logic;

    signal FIN_ANDGate_214, RDY_ANDGate_214 : std_logic;

    signal FIN_ANDGate_215, RDY_ANDGate_215 : std_logic;

    signal FIN_ANDGate_216, RDY_ANDGate_216 : std_logic;

    signal FIN_ANDGate_217, RDY_ANDGate_217 : std_logic;

    signal FIN_ANDGate_218, RDY_ANDGate_218 : std_logic;

    signal FIN_ANDGate_219, RDY_ANDGate_219 : std_logic;

    signal FIN_ANDGate_220, RDY_ANDGate_220 : std_logic;

    signal FIN_ANDGate_221, RDY_ANDGate_221 : std_logic;

    signal FIN_ANDGate_222, RDY_ANDGate_222 : std_logic;

    signal FIN_ANDGate_223, RDY_ANDGate_223 : std_logic;

    signal FIN_ANDGate_224, RDY_ANDGate_224 : std_logic;

    signal FIN_ANDGate_225, RDY_ANDGate_225 : std_logic;

    signal FIN_ANDGate_226, RDY_ANDGate_226 : std_logic;

    signal FIN_ANDGate_227, RDY_ANDGate_227 : std_logic;

    signal FIN_ANDGate_228, RDY_ANDGate_228 : std_logic;

    signal FIN_ANDGate_229, RDY_ANDGate_229 : std_logic;

    signal FIN_ANDGate_230, RDY_ANDGate_230 : std_logic;

    signal FIN_ANDGate_231, RDY_ANDGate_231 : std_logic;

    signal FIN_ANDGate_232, RDY_ANDGate_232 : std_logic;

    signal FIN_ANDGate_233, RDY_ANDGate_233 : std_logic;

    signal FIN_ANDGate_234, RDY_ANDGate_234 : std_logic;

    signal FIN_ANDGate_235, RDY_ANDGate_235 : std_logic;

    signal FIN_ANDGate_236, RDY_ANDGate_236 : std_logic;

    signal FIN_ANDGate_237, RDY_ANDGate_237 : std_logic;

    signal FIN_ANDGate_238, RDY_ANDGate_238 : std_logic;

    signal FIN_ANDGate_239, RDY_ANDGate_239 : std_logic;

    signal FIN_ANDGate_240, RDY_ANDGate_240 : std_logic;

    signal FIN_ANDGate_241, RDY_ANDGate_241 : std_logic;

    signal FIN_ANDGate_242, RDY_ANDGate_242 : std_logic;

    signal FIN_ANDGate_243, RDY_ANDGate_243 : std_logic;

    signal FIN_ANDGate_244, RDY_ANDGate_244 : std_logic;

    signal FIN_ANDGate_245, RDY_ANDGate_245 : std_logic;

    signal FIN_ANDGate_246, RDY_ANDGate_246 : std_logic;

    signal FIN_ANDGate_247, RDY_ANDGate_247 : std_logic;

    signal FIN_ANDGate_248, RDY_ANDGate_248 : std_logic;

    signal FIN_ANDGate_249, RDY_ANDGate_249 : std_logic;

    signal FIN_ANDGate_250, RDY_ANDGate_250 : std_logic;

    signal FIN_ANDGate_251, RDY_ANDGate_251 : std_logic;

    signal FIN_ANDGate_252, RDY_ANDGate_252 : std_logic;

    signal FIN_ANDGate_253, RDY_ANDGate_253 : std_logic;

    signal FIN_ANDGate_254, RDY_ANDGate_254 : std_logic;

    signal FIN_ANDGate_255, RDY_ANDGate_255 : std_logic;


    -- The primary ready driver signal
    signal RDY : std_logic;

begin


    -- Entity  NOTGate_0 signals
    NOTGate_0: entity work.NOTGate_0
    port map (
        -- Input bus DecoderInput_0
        m_input_Value => DecoderInput_0_Value,


        -- Output bus DecoderNOTInput_0
        output_0_Value => DecoderNOTInput_0_Value,



        CLK => CLK,
        RDY => RDY_NOTGate_0,
        FIN => FIN_NOTGate_0,
        ENB => ENB,
        RST => RST
    );


    -- Entity  NOTGate_1 signals
    NOTGate_1: entity work.NOTGate_1
    port map (
        -- Input bus DecoderInput_1
        m_input_Value => DecoderInput_1_Value,


        -- Output bus DecoderNOTInput_1
        output_1_Value => DecoderNOTInput_1_Value,



        CLK => CLK,
        RDY => RDY_NOTGate_1,
        FIN => FIN_NOTGate_1,
        ENB => ENB,
        RST => RST
    );


    -- Entity  NOTGate_2 signals
    NOTGate_2: entity work.NOTGate_2
    port map (
        -- Input bus DecoderInput_2
        m_input_Value => DecoderInput_2_Value,


        -- Output bus DecoderNOTInput_2
        output_2_Value => DecoderNOTInput_2_Value,



        CLK => CLK,
        RDY => RDY_NOTGate_2,
        FIN => FIN_NOTGate_2,
        ENB => ENB,
        RST => RST
    );


    -- Entity  NOTGate_3 signals
    NOTGate_3: entity work.NOTGate_3
    port map (
        -- Input bus DecoderInput_3
        m_input_Value => DecoderInput_3_Value,


        -- Output bus DecoderNOTInput_3
        output_3_Value => DecoderNOTInput_3_Value,



        CLK => CLK,
        RDY => RDY_NOTGate_3,
        FIN => FIN_NOTGate_3,
        ENB => ENB,
        RST => RST
    );


    -- Entity  NOTGate_4 signals
    NOTGate_4: entity work.NOTGate_4
    port map (
        -- Input bus DecoderInput_4
        m_input_Value => DecoderInput_4_Value,


        -- Output bus DecoderNOTInput_4
        output_4_Value => DecoderNOTInput_4_Value,



        CLK => CLK,
        RDY => RDY_NOTGate_4,
        FIN => FIN_NOTGate_4,
        ENB => ENB,
        RST => RST
    );


    -- Entity  NOTGate_5 signals
    NOTGate_5: entity work.NOTGate_5
    port map (
        -- Input bus DecoderInput_5
        m_input_Value => DecoderInput_5_Value,


        -- Output bus DecoderNOTInput_5
        output_5_Value => DecoderNOTInput_5_Value,



        CLK => CLK,
        RDY => RDY_NOTGate_5,
        FIN => FIN_NOTGate_5,
        ENB => ENB,
        RST => RST
    );


    -- Entity  NOTGate_6 signals
    NOTGate_6: entity work.NOTGate_6
    port map (
        -- Input bus DecoderInput_6
        m_input_Value => DecoderInput_6_Value,


        -- Output bus DecoderNOTInput_6
        output_6_Value => DecoderNOTInput_6_Value,



        CLK => CLK,
        RDY => RDY_NOTGate_6,
        FIN => FIN_NOTGate_6,
        ENB => ENB,
        RST => RST
    );


    -- Entity  NOTGate_7 signals
    NOTGate_7: entity work.NOTGate_7
    port map (
        -- Input bus DecoderInput_7
        m_input_Value => DecoderInput_7_Value,


        -- Output bus DecoderNOTInput_7
        output_7_Value => DecoderNOTInput_7_Value,



        CLK => CLK,
        RDY => RDY_NOTGate_7,
        FIN => FIN_NOTGate_7,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_0 signals
    ANDGate_0: entity work.ANDGate_0
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_0
        output_0_Value => DecoderOutput_0_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_0,
        FIN => FIN_ANDGate_0,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_1 signals
    ANDGate_1: entity work.ANDGate_1
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_1
        output_1_Value => DecoderOutput_1_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_1,
        FIN => FIN_ANDGate_1,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_2 signals
    ANDGate_2: entity work.ANDGate_2
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_2
        output_2_Value => DecoderOutput_2_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_2,
        FIN => FIN_ANDGate_2,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_3 signals
    ANDGate_3: entity work.ANDGate_3
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_3
        output_3_Value => DecoderOutput_3_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_3,
        FIN => FIN_ANDGate_3,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_4 signals
    ANDGate_4: entity work.ANDGate_4
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_4
        output_4_Value => DecoderOutput_4_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_4,
        FIN => FIN_ANDGate_4,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_5 signals
    ANDGate_5: entity work.ANDGate_5
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_5
        output_5_Value => DecoderOutput_5_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_5,
        FIN => FIN_ANDGate_5,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_6 signals
    ANDGate_6: entity work.ANDGate_6
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_6
        output_6_Value => DecoderOutput_6_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_6,
        FIN => FIN_ANDGate_6,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_7 signals
    ANDGate_7: entity work.ANDGate_7
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_7
        output_7_Value => DecoderOutput_7_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_7,
        FIN => FIN_ANDGate_7,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_8 signals
    ANDGate_8: entity work.ANDGate_8
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_8
        output_8_Value => DecoderOutput_8_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_8,
        FIN => FIN_ANDGate_8,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_9 signals
    ANDGate_9: entity work.ANDGate_9
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_9
        output_9_Value => DecoderOutput_9_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_9,
        FIN => FIN_ANDGate_9,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_10 signals
    ANDGate_10: entity work.ANDGate_10
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_10
        output_10_Value => DecoderOutput_10_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_10,
        FIN => FIN_ANDGate_10,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_11 signals
    ANDGate_11: entity work.ANDGate_11
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_11
        output_11_Value => DecoderOutput_11_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_11,
        FIN => FIN_ANDGate_11,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_12 signals
    ANDGate_12: entity work.ANDGate_12
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_12
        output_12_Value => DecoderOutput_12_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_12,
        FIN => FIN_ANDGate_12,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_13 signals
    ANDGate_13: entity work.ANDGate_13
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_13
        output_13_Value => DecoderOutput_13_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_13,
        FIN => FIN_ANDGate_13,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_14 signals
    ANDGate_14: entity work.ANDGate_14
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_14
        output_14_Value => DecoderOutput_14_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_14,
        FIN => FIN_ANDGate_14,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_15 signals
    ANDGate_15: entity work.ANDGate_15
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_15
        output_15_Value => DecoderOutput_15_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_15,
        FIN => FIN_ANDGate_15,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_16 signals
    ANDGate_16: entity work.ANDGate_16
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_16
        output_16_Value => DecoderOutput_16_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_16,
        FIN => FIN_ANDGate_16,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_17 signals
    ANDGate_17: entity work.ANDGate_17
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_17
        output_17_Value => DecoderOutput_17_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_17,
        FIN => FIN_ANDGate_17,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_18 signals
    ANDGate_18: entity work.ANDGate_18
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_18
        output_18_Value => DecoderOutput_18_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_18,
        FIN => FIN_ANDGate_18,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_19 signals
    ANDGate_19: entity work.ANDGate_19
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_19
        output_19_Value => DecoderOutput_19_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_19,
        FIN => FIN_ANDGate_19,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_20 signals
    ANDGate_20: entity work.ANDGate_20
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_20
        output_20_Value => DecoderOutput_20_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_20,
        FIN => FIN_ANDGate_20,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_21 signals
    ANDGate_21: entity work.ANDGate_21
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_21
        output_21_Value => DecoderOutput_21_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_21,
        FIN => FIN_ANDGate_21,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_22 signals
    ANDGate_22: entity work.ANDGate_22
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_22
        output_22_Value => DecoderOutput_22_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_22,
        FIN => FIN_ANDGate_22,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_23 signals
    ANDGate_23: entity work.ANDGate_23
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_23
        output_23_Value => DecoderOutput_23_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_23,
        FIN => FIN_ANDGate_23,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_24 signals
    ANDGate_24: entity work.ANDGate_24
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_24
        output_24_Value => DecoderOutput_24_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_24,
        FIN => FIN_ANDGate_24,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_25 signals
    ANDGate_25: entity work.ANDGate_25
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_25
        output_25_Value => DecoderOutput_25_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_25,
        FIN => FIN_ANDGate_25,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_26 signals
    ANDGate_26: entity work.ANDGate_26
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_26
        output_26_Value => DecoderOutput_26_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_26,
        FIN => FIN_ANDGate_26,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_27 signals
    ANDGate_27: entity work.ANDGate_27
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_27
        output_27_Value => DecoderOutput_27_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_27,
        FIN => FIN_ANDGate_27,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_28 signals
    ANDGate_28: entity work.ANDGate_28
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_28
        output_28_Value => DecoderOutput_28_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_28,
        FIN => FIN_ANDGate_28,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_29 signals
    ANDGate_29: entity work.ANDGate_29
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_29
        output_29_Value => DecoderOutput_29_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_29,
        FIN => FIN_ANDGate_29,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_30 signals
    ANDGate_30: entity work.ANDGate_30
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_30
        output_30_Value => DecoderOutput_30_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_30,
        FIN => FIN_ANDGate_30,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_31 signals
    ANDGate_31: entity work.ANDGate_31
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_31
        output_31_Value => DecoderOutput_31_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_31,
        FIN => FIN_ANDGate_31,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_32 signals
    ANDGate_32: entity work.ANDGate_32
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_32
        output_32_Value => DecoderOutput_32_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_32,
        FIN => FIN_ANDGate_32,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_33 signals
    ANDGate_33: entity work.ANDGate_33
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_33
        output_33_Value => DecoderOutput_33_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_33,
        FIN => FIN_ANDGate_33,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_34 signals
    ANDGate_34: entity work.ANDGate_34
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_34
        output_34_Value => DecoderOutput_34_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_34,
        FIN => FIN_ANDGate_34,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_35 signals
    ANDGate_35: entity work.ANDGate_35
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_35
        output_35_Value => DecoderOutput_35_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_35,
        FIN => FIN_ANDGate_35,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_36 signals
    ANDGate_36: entity work.ANDGate_36
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_36
        output_36_Value => DecoderOutput_36_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_36,
        FIN => FIN_ANDGate_36,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_37 signals
    ANDGate_37: entity work.ANDGate_37
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_37
        output_37_Value => DecoderOutput_37_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_37,
        FIN => FIN_ANDGate_37,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_38 signals
    ANDGate_38: entity work.ANDGate_38
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_38
        output_38_Value => DecoderOutput_38_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_38,
        FIN => FIN_ANDGate_38,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_39 signals
    ANDGate_39: entity work.ANDGate_39
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_39
        output_39_Value => DecoderOutput_39_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_39,
        FIN => FIN_ANDGate_39,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_40 signals
    ANDGate_40: entity work.ANDGate_40
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_40
        output_40_Value => DecoderOutput_40_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_40,
        FIN => FIN_ANDGate_40,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_41 signals
    ANDGate_41: entity work.ANDGate_41
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_41
        output_41_Value => DecoderOutput_41_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_41,
        FIN => FIN_ANDGate_41,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_42 signals
    ANDGate_42: entity work.ANDGate_42
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_42
        output_42_Value => DecoderOutput_42_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_42,
        FIN => FIN_ANDGate_42,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_43 signals
    ANDGate_43: entity work.ANDGate_43
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_43
        output_43_Value => DecoderOutput_43_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_43,
        FIN => FIN_ANDGate_43,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_44 signals
    ANDGate_44: entity work.ANDGate_44
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_44
        output_44_Value => DecoderOutput_44_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_44,
        FIN => FIN_ANDGate_44,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_45 signals
    ANDGate_45: entity work.ANDGate_45
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_45
        output_45_Value => DecoderOutput_45_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_45,
        FIN => FIN_ANDGate_45,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_46 signals
    ANDGate_46: entity work.ANDGate_46
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_46
        output_46_Value => DecoderOutput_46_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_46,
        FIN => FIN_ANDGate_46,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_47 signals
    ANDGate_47: entity work.ANDGate_47
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_47
        output_47_Value => DecoderOutput_47_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_47,
        FIN => FIN_ANDGate_47,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_48 signals
    ANDGate_48: entity work.ANDGate_48
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_48
        output_48_Value => DecoderOutput_48_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_48,
        FIN => FIN_ANDGate_48,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_49 signals
    ANDGate_49: entity work.ANDGate_49
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_49
        output_49_Value => DecoderOutput_49_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_49,
        FIN => FIN_ANDGate_49,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_50 signals
    ANDGate_50: entity work.ANDGate_50
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_50
        output_50_Value => DecoderOutput_50_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_50,
        FIN => FIN_ANDGate_50,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_51 signals
    ANDGate_51: entity work.ANDGate_51
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_51
        output_51_Value => DecoderOutput_51_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_51,
        FIN => FIN_ANDGate_51,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_52 signals
    ANDGate_52: entity work.ANDGate_52
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_52
        output_52_Value => DecoderOutput_52_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_52,
        FIN => FIN_ANDGate_52,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_53 signals
    ANDGate_53: entity work.ANDGate_53
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_53
        output_53_Value => DecoderOutput_53_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_53,
        FIN => FIN_ANDGate_53,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_54 signals
    ANDGate_54: entity work.ANDGate_54
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_54
        output_54_Value => DecoderOutput_54_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_54,
        FIN => FIN_ANDGate_54,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_55 signals
    ANDGate_55: entity work.ANDGate_55
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_55
        output_55_Value => DecoderOutput_55_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_55,
        FIN => FIN_ANDGate_55,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_56 signals
    ANDGate_56: entity work.ANDGate_56
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_56
        output_56_Value => DecoderOutput_56_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_56,
        FIN => FIN_ANDGate_56,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_57 signals
    ANDGate_57: entity work.ANDGate_57
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_57
        output_57_Value => DecoderOutput_57_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_57,
        FIN => FIN_ANDGate_57,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_58 signals
    ANDGate_58: entity work.ANDGate_58
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_58
        output_58_Value => DecoderOutput_58_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_58,
        FIN => FIN_ANDGate_58,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_59 signals
    ANDGate_59: entity work.ANDGate_59
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_59
        output_59_Value => DecoderOutput_59_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_59,
        FIN => FIN_ANDGate_59,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_60 signals
    ANDGate_60: entity work.ANDGate_60
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_60
        output_60_Value => DecoderOutput_60_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_60,
        FIN => FIN_ANDGate_60,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_61 signals
    ANDGate_61: entity work.ANDGate_61
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_61
        output_61_Value => DecoderOutput_61_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_61,
        FIN => FIN_ANDGate_61,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_62 signals
    ANDGate_62: entity work.ANDGate_62
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_62
        output_62_Value => DecoderOutput_62_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_62,
        FIN => FIN_ANDGate_62,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_63 signals
    ANDGate_63: entity work.ANDGate_63
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_63
        output_63_Value => DecoderOutput_63_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_63,
        FIN => FIN_ANDGate_63,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_64 signals
    ANDGate_64: entity work.ANDGate_64
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_64
        output_64_Value => DecoderOutput_64_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_64,
        FIN => FIN_ANDGate_64,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_65 signals
    ANDGate_65: entity work.ANDGate_65
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_65
        output_65_Value => DecoderOutput_65_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_65,
        FIN => FIN_ANDGate_65,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_66 signals
    ANDGate_66: entity work.ANDGate_66
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_66
        output_66_Value => DecoderOutput_66_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_66,
        FIN => FIN_ANDGate_66,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_67 signals
    ANDGate_67: entity work.ANDGate_67
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_67
        output_67_Value => DecoderOutput_67_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_67,
        FIN => FIN_ANDGate_67,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_68 signals
    ANDGate_68: entity work.ANDGate_68
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_68
        output_68_Value => DecoderOutput_68_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_68,
        FIN => FIN_ANDGate_68,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_69 signals
    ANDGate_69: entity work.ANDGate_69
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_69
        output_69_Value => DecoderOutput_69_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_69,
        FIN => FIN_ANDGate_69,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_70 signals
    ANDGate_70: entity work.ANDGate_70
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_70
        output_70_Value => DecoderOutput_70_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_70,
        FIN => FIN_ANDGate_70,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_71 signals
    ANDGate_71: entity work.ANDGate_71
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_71
        output_71_Value => DecoderOutput_71_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_71,
        FIN => FIN_ANDGate_71,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_72 signals
    ANDGate_72: entity work.ANDGate_72
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_72
        output_72_Value => DecoderOutput_72_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_72,
        FIN => FIN_ANDGate_72,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_73 signals
    ANDGate_73: entity work.ANDGate_73
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_73
        output_73_Value => DecoderOutput_73_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_73,
        FIN => FIN_ANDGate_73,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_74 signals
    ANDGate_74: entity work.ANDGate_74
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_74
        output_74_Value => DecoderOutput_74_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_74,
        FIN => FIN_ANDGate_74,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_75 signals
    ANDGate_75: entity work.ANDGate_75
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_75
        output_75_Value => DecoderOutput_75_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_75,
        FIN => FIN_ANDGate_75,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_76 signals
    ANDGate_76: entity work.ANDGate_76
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_76
        output_76_Value => DecoderOutput_76_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_76,
        FIN => FIN_ANDGate_76,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_77 signals
    ANDGate_77: entity work.ANDGate_77
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_77
        output_77_Value => DecoderOutput_77_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_77,
        FIN => FIN_ANDGate_77,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_78 signals
    ANDGate_78: entity work.ANDGate_78
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_78
        output_78_Value => DecoderOutput_78_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_78,
        FIN => FIN_ANDGate_78,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_79 signals
    ANDGate_79: entity work.ANDGate_79
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_79
        output_79_Value => DecoderOutput_79_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_79,
        FIN => FIN_ANDGate_79,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_80 signals
    ANDGate_80: entity work.ANDGate_80
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_80
        output_80_Value => DecoderOutput_80_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_80,
        FIN => FIN_ANDGate_80,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_81 signals
    ANDGate_81: entity work.ANDGate_81
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_81
        output_81_Value => DecoderOutput_81_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_81,
        FIN => FIN_ANDGate_81,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_82 signals
    ANDGate_82: entity work.ANDGate_82
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_82
        output_82_Value => DecoderOutput_82_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_82,
        FIN => FIN_ANDGate_82,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_83 signals
    ANDGate_83: entity work.ANDGate_83
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_83
        output_83_Value => DecoderOutput_83_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_83,
        FIN => FIN_ANDGate_83,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_84 signals
    ANDGate_84: entity work.ANDGate_84
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_84
        output_84_Value => DecoderOutput_84_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_84,
        FIN => FIN_ANDGate_84,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_85 signals
    ANDGate_85: entity work.ANDGate_85
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_85
        output_85_Value => DecoderOutput_85_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_85,
        FIN => FIN_ANDGate_85,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_86 signals
    ANDGate_86: entity work.ANDGate_86
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_86
        output_86_Value => DecoderOutput_86_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_86,
        FIN => FIN_ANDGate_86,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_87 signals
    ANDGate_87: entity work.ANDGate_87
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_87
        output_87_Value => DecoderOutput_87_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_87,
        FIN => FIN_ANDGate_87,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_88 signals
    ANDGate_88: entity work.ANDGate_88
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_88
        output_88_Value => DecoderOutput_88_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_88,
        FIN => FIN_ANDGate_88,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_89 signals
    ANDGate_89: entity work.ANDGate_89
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_89
        output_89_Value => DecoderOutput_89_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_89,
        FIN => FIN_ANDGate_89,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_90 signals
    ANDGate_90: entity work.ANDGate_90
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_90
        output_90_Value => DecoderOutput_90_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_90,
        FIN => FIN_ANDGate_90,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_91 signals
    ANDGate_91: entity work.ANDGate_91
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_91
        output_91_Value => DecoderOutput_91_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_91,
        FIN => FIN_ANDGate_91,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_92 signals
    ANDGate_92: entity work.ANDGate_92
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_92
        output_92_Value => DecoderOutput_92_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_92,
        FIN => FIN_ANDGate_92,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_93 signals
    ANDGate_93: entity work.ANDGate_93
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_93
        output_93_Value => DecoderOutput_93_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_93,
        FIN => FIN_ANDGate_93,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_94 signals
    ANDGate_94: entity work.ANDGate_94
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_94
        output_94_Value => DecoderOutput_94_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_94,
        FIN => FIN_ANDGate_94,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_95 signals
    ANDGate_95: entity work.ANDGate_95
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_95
        output_95_Value => DecoderOutput_95_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_95,
        FIN => FIN_ANDGate_95,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_96 signals
    ANDGate_96: entity work.ANDGate_96
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_96
        output_96_Value => DecoderOutput_96_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_96,
        FIN => FIN_ANDGate_96,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_97 signals
    ANDGate_97: entity work.ANDGate_97
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_97
        output_97_Value => DecoderOutput_97_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_97,
        FIN => FIN_ANDGate_97,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_98 signals
    ANDGate_98: entity work.ANDGate_98
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_98
        output_98_Value => DecoderOutput_98_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_98,
        FIN => FIN_ANDGate_98,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_99 signals
    ANDGate_99: entity work.ANDGate_99
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_99
        output_99_Value => DecoderOutput_99_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_99,
        FIN => FIN_ANDGate_99,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_100 signals
    ANDGate_100: entity work.ANDGate_100
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_100
        output_100_Value => DecoderOutput_100_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_100,
        FIN => FIN_ANDGate_100,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_101 signals
    ANDGate_101: entity work.ANDGate_101
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_101
        output_101_Value => DecoderOutput_101_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_101,
        FIN => FIN_ANDGate_101,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_102 signals
    ANDGate_102: entity work.ANDGate_102
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_102
        output_102_Value => DecoderOutput_102_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_102,
        FIN => FIN_ANDGate_102,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_103 signals
    ANDGate_103: entity work.ANDGate_103
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_103
        output_103_Value => DecoderOutput_103_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_103,
        FIN => FIN_ANDGate_103,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_104 signals
    ANDGate_104: entity work.ANDGate_104
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_104
        output_104_Value => DecoderOutput_104_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_104,
        FIN => FIN_ANDGate_104,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_105 signals
    ANDGate_105: entity work.ANDGate_105
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_105
        output_105_Value => DecoderOutput_105_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_105,
        FIN => FIN_ANDGate_105,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_106 signals
    ANDGate_106: entity work.ANDGate_106
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_106
        output_106_Value => DecoderOutput_106_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_106,
        FIN => FIN_ANDGate_106,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_107 signals
    ANDGate_107: entity work.ANDGate_107
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_107
        output_107_Value => DecoderOutput_107_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_107,
        FIN => FIN_ANDGate_107,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_108 signals
    ANDGate_108: entity work.ANDGate_108
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_108
        output_108_Value => DecoderOutput_108_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_108,
        FIN => FIN_ANDGate_108,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_109 signals
    ANDGate_109: entity work.ANDGate_109
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_109
        output_109_Value => DecoderOutput_109_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_109,
        FIN => FIN_ANDGate_109,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_110 signals
    ANDGate_110: entity work.ANDGate_110
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_110
        output_110_Value => DecoderOutput_110_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_110,
        FIN => FIN_ANDGate_110,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_111 signals
    ANDGate_111: entity work.ANDGate_111
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_111
        output_111_Value => DecoderOutput_111_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_111,
        FIN => FIN_ANDGate_111,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_112 signals
    ANDGate_112: entity work.ANDGate_112
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_112
        output_112_Value => DecoderOutput_112_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_112,
        FIN => FIN_ANDGate_112,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_113 signals
    ANDGate_113: entity work.ANDGate_113
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_113
        output_113_Value => DecoderOutput_113_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_113,
        FIN => FIN_ANDGate_113,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_114 signals
    ANDGate_114: entity work.ANDGate_114
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_114
        output_114_Value => DecoderOutput_114_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_114,
        FIN => FIN_ANDGate_114,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_115 signals
    ANDGate_115: entity work.ANDGate_115
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_115
        output_115_Value => DecoderOutput_115_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_115,
        FIN => FIN_ANDGate_115,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_116 signals
    ANDGate_116: entity work.ANDGate_116
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_116
        output_116_Value => DecoderOutput_116_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_116,
        FIN => FIN_ANDGate_116,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_117 signals
    ANDGate_117: entity work.ANDGate_117
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_117
        output_117_Value => DecoderOutput_117_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_117,
        FIN => FIN_ANDGate_117,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_118 signals
    ANDGate_118: entity work.ANDGate_118
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_118
        output_118_Value => DecoderOutput_118_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_118,
        FIN => FIN_ANDGate_118,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_119 signals
    ANDGate_119: entity work.ANDGate_119
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_119
        output_119_Value => DecoderOutput_119_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_119,
        FIN => FIN_ANDGate_119,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_120 signals
    ANDGate_120: entity work.ANDGate_120
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_120
        output_120_Value => DecoderOutput_120_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_120,
        FIN => FIN_ANDGate_120,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_121 signals
    ANDGate_121: entity work.ANDGate_121
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_121
        output_121_Value => DecoderOutput_121_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_121,
        FIN => FIN_ANDGate_121,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_122 signals
    ANDGate_122: entity work.ANDGate_122
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_122
        output_122_Value => DecoderOutput_122_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_122,
        FIN => FIN_ANDGate_122,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_123 signals
    ANDGate_123: entity work.ANDGate_123
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_123
        output_123_Value => DecoderOutput_123_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_123,
        FIN => FIN_ANDGate_123,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_124 signals
    ANDGate_124: entity work.ANDGate_124
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_124
        output_124_Value => DecoderOutput_124_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_124,
        FIN => FIN_ANDGate_124,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_125 signals
    ANDGate_125: entity work.ANDGate_125
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_125
        output_125_Value => DecoderOutput_125_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_125,
        FIN => FIN_ANDGate_125,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_126 signals
    ANDGate_126: entity work.ANDGate_126
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_126
        output_126_Value => DecoderOutput_126_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_126,
        FIN => FIN_ANDGate_126,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_127 signals
    ANDGate_127: entity work.ANDGate_127
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderNOTInput_7
        m_input_NOT_7_Value => DecoderNOTInput_7_Value,


        -- Output bus DecoderOutput_127
        output_127_Value => DecoderOutput_127_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_127,
        FIN => FIN_ANDGate_127,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_128 signals
    ANDGate_128: entity work.ANDGate_128
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_128
        output_128_Value => DecoderOutput_128_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_128,
        FIN => FIN_ANDGate_128,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_129 signals
    ANDGate_129: entity work.ANDGate_129
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_129
        output_129_Value => DecoderOutput_129_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_129,
        FIN => FIN_ANDGate_129,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_130 signals
    ANDGate_130: entity work.ANDGate_130
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_130
        output_130_Value => DecoderOutput_130_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_130,
        FIN => FIN_ANDGate_130,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_131 signals
    ANDGate_131: entity work.ANDGate_131
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_131
        output_131_Value => DecoderOutput_131_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_131,
        FIN => FIN_ANDGate_131,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_132 signals
    ANDGate_132: entity work.ANDGate_132
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_132
        output_132_Value => DecoderOutput_132_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_132,
        FIN => FIN_ANDGate_132,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_133 signals
    ANDGate_133: entity work.ANDGate_133
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_133
        output_133_Value => DecoderOutput_133_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_133,
        FIN => FIN_ANDGate_133,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_134 signals
    ANDGate_134: entity work.ANDGate_134
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_134
        output_134_Value => DecoderOutput_134_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_134,
        FIN => FIN_ANDGate_134,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_135 signals
    ANDGate_135: entity work.ANDGate_135
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_135
        output_135_Value => DecoderOutput_135_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_135,
        FIN => FIN_ANDGate_135,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_136 signals
    ANDGate_136: entity work.ANDGate_136
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_136
        output_136_Value => DecoderOutput_136_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_136,
        FIN => FIN_ANDGate_136,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_137 signals
    ANDGate_137: entity work.ANDGate_137
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_137
        output_137_Value => DecoderOutput_137_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_137,
        FIN => FIN_ANDGate_137,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_138 signals
    ANDGate_138: entity work.ANDGate_138
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_138
        output_138_Value => DecoderOutput_138_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_138,
        FIN => FIN_ANDGate_138,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_139 signals
    ANDGate_139: entity work.ANDGate_139
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_139
        output_139_Value => DecoderOutput_139_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_139,
        FIN => FIN_ANDGate_139,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_140 signals
    ANDGate_140: entity work.ANDGate_140
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_140
        output_140_Value => DecoderOutput_140_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_140,
        FIN => FIN_ANDGate_140,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_141 signals
    ANDGate_141: entity work.ANDGate_141
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_141
        output_141_Value => DecoderOutput_141_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_141,
        FIN => FIN_ANDGate_141,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_142 signals
    ANDGate_142: entity work.ANDGate_142
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_142
        output_142_Value => DecoderOutput_142_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_142,
        FIN => FIN_ANDGate_142,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_143 signals
    ANDGate_143: entity work.ANDGate_143
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_143
        output_143_Value => DecoderOutput_143_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_143,
        FIN => FIN_ANDGate_143,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_144 signals
    ANDGate_144: entity work.ANDGate_144
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_144
        output_144_Value => DecoderOutput_144_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_144,
        FIN => FIN_ANDGate_144,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_145 signals
    ANDGate_145: entity work.ANDGate_145
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_145
        output_145_Value => DecoderOutput_145_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_145,
        FIN => FIN_ANDGate_145,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_146 signals
    ANDGate_146: entity work.ANDGate_146
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_146
        output_146_Value => DecoderOutput_146_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_146,
        FIN => FIN_ANDGate_146,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_147 signals
    ANDGate_147: entity work.ANDGate_147
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_147
        output_147_Value => DecoderOutput_147_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_147,
        FIN => FIN_ANDGate_147,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_148 signals
    ANDGate_148: entity work.ANDGate_148
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_148
        output_148_Value => DecoderOutput_148_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_148,
        FIN => FIN_ANDGate_148,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_149 signals
    ANDGate_149: entity work.ANDGate_149
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_149
        output_149_Value => DecoderOutput_149_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_149,
        FIN => FIN_ANDGate_149,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_150 signals
    ANDGate_150: entity work.ANDGate_150
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_150
        output_150_Value => DecoderOutput_150_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_150,
        FIN => FIN_ANDGate_150,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_151 signals
    ANDGate_151: entity work.ANDGate_151
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_151
        output_151_Value => DecoderOutput_151_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_151,
        FIN => FIN_ANDGate_151,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_152 signals
    ANDGate_152: entity work.ANDGate_152
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_152
        output_152_Value => DecoderOutput_152_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_152,
        FIN => FIN_ANDGate_152,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_153 signals
    ANDGate_153: entity work.ANDGate_153
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_153
        output_153_Value => DecoderOutput_153_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_153,
        FIN => FIN_ANDGate_153,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_154 signals
    ANDGate_154: entity work.ANDGate_154
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_154
        output_154_Value => DecoderOutput_154_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_154,
        FIN => FIN_ANDGate_154,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_155 signals
    ANDGate_155: entity work.ANDGate_155
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_155
        output_155_Value => DecoderOutput_155_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_155,
        FIN => FIN_ANDGate_155,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_156 signals
    ANDGate_156: entity work.ANDGate_156
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_156
        output_156_Value => DecoderOutput_156_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_156,
        FIN => FIN_ANDGate_156,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_157 signals
    ANDGate_157: entity work.ANDGate_157
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_157
        output_157_Value => DecoderOutput_157_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_157,
        FIN => FIN_ANDGate_157,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_158 signals
    ANDGate_158: entity work.ANDGate_158
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_158
        output_158_Value => DecoderOutput_158_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_158,
        FIN => FIN_ANDGate_158,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_159 signals
    ANDGate_159: entity work.ANDGate_159
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_159
        output_159_Value => DecoderOutput_159_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_159,
        FIN => FIN_ANDGate_159,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_160 signals
    ANDGate_160: entity work.ANDGate_160
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_160
        output_160_Value => DecoderOutput_160_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_160,
        FIN => FIN_ANDGate_160,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_161 signals
    ANDGate_161: entity work.ANDGate_161
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_161
        output_161_Value => DecoderOutput_161_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_161,
        FIN => FIN_ANDGate_161,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_162 signals
    ANDGate_162: entity work.ANDGate_162
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_162
        output_162_Value => DecoderOutput_162_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_162,
        FIN => FIN_ANDGate_162,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_163 signals
    ANDGate_163: entity work.ANDGate_163
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_163
        output_163_Value => DecoderOutput_163_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_163,
        FIN => FIN_ANDGate_163,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_164 signals
    ANDGate_164: entity work.ANDGate_164
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_164
        output_164_Value => DecoderOutput_164_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_164,
        FIN => FIN_ANDGate_164,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_165 signals
    ANDGate_165: entity work.ANDGate_165
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_165
        output_165_Value => DecoderOutput_165_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_165,
        FIN => FIN_ANDGate_165,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_166 signals
    ANDGate_166: entity work.ANDGate_166
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_166
        output_166_Value => DecoderOutput_166_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_166,
        FIN => FIN_ANDGate_166,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_167 signals
    ANDGate_167: entity work.ANDGate_167
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_167
        output_167_Value => DecoderOutput_167_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_167,
        FIN => FIN_ANDGate_167,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_168 signals
    ANDGate_168: entity work.ANDGate_168
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_168
        output_168_Value => DecoderOutput_168_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_168,
        FIN => FIN_ANDGate_168,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_169 signals
    ANDGate_169: entity work.ANDGate_169
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_169
        output_169_Value => DecoderOutput_169_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_169,
        FIN => FIN_ANDGate_169,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_170 signals
    ANDGate_170: entity work.ANDGate_170
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_170
        output_170_Value => DecoderOutput_170_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_170,
        FIN => FIN_ANDGate_170,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_171 signals
    ANDGate_171: entity work.ANDGate_171
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_171
        output_171_Value => DecoderOutput_171_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_171,
        FIN => FIN_ANDGate_171,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_172 signals
    ANDGate_172: entity work.ANDGate_172
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_172
        output_172_Value => DecoderOutput_172_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_172,
        FIN => FIN_ANDGate_172,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_173 signals
    ANDGate_173: entity work.ANDGate_173
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_173
        output_173_Value => DecoderOutput_173_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_173,
        FIN => FIN_ANDGate_173,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_174 signals
    ANDGate_174: entity work.ANDGate_174
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_174
        output_174_Value => DecoderOutput_174_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_174,
        FIN => FIN_ANDGate_174,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_175 signals
    ANDGate_175: entity work.ANDGate_175
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_175
        output_175_Value => DecoderOutput_175_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_175,
        FIN => FIN_ANDGate_175,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_176 signals
    ANDGate_176: entity work.ANDGate_176
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_176
        output_176_Value => DecoderOutput_176_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_176,
        FIN => FIN_ANDGate_176,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_177 signals
    ANDGate_177: entity work.ANDGate_177
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_177
        output_177_Value => DecoderOutput_177_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_177,
        FIN => FIN_ANDGate_177,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_178 signals
    ANDGate_178: entity work.ANDGate_178
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_178
        output_178_Value => DecoderOutput_178_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_178,
        FIN => FIN_ANDGate_178,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_179 signals
    ANDGate_179: entity work.ANDGate_179
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_179
        output_179_Value => DecoderOutput_179_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_179,
        FIN => FIN_ANDGate_179,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_180 signals
    ANDGate_180: entity work.ANDGate_180
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_180
        output_180_Value => DecoderOutput_180_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_180,
        FIN => FIN_ANDGate_180,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_181 signals
    ANDGate_181: entity work.ANDGate_181
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_181
        output_181_Value => DecoderOutput_181_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_181,
        FIN => FIN_ANDGate_181,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_182 signals
    ANDGate_182: entity work.ANDGate_182
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_182
        output_182_Value => DecoderOutput_182_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_182,
        FIN => FIN_ANDGate_182,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_183 signals
    ANDGate_183: entity work.ANDGate_183
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_183
        output_183_Value => DecoderOutput_183_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_183,
        FIN => FIN_ANDGate_183,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_184 signals
    ANDGate_184: entity work.ANDGate_184
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_184
        output_184_Value => DecoderOutput_184_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_184,
        FIN => FIN_ANDGate_184,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_185 signals
    ANDGate_185: entity work.ANDGate_185
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_185
        output_185_Value => DecoderOutput_185_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_185,
        FIN => FIN_ANDGate_185,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_186 signals
    ANDGate_186: entity work.ANDGate_186
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_186
        output_186_Value => DecoderOutput_186_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_186,
        FIN => FIN_ANDGate_186,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_187 signals
    ANDGate_187: entity work.ANDGate_187
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_187
        output_187_Value => DecoderOutput_187_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_187,
        FIN => FIN_ANDGate_187,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_188 signals
    ANDGate_188: entity work.ANDGate_188
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_188
        output_188_Value => DecoderOutput_188_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_188,
        FIN => FIN_ANDGate_188,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_189 signals
    ANDGate_189: entity work.ANDGate_189
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_189
        output_189_Value => DecoderOutput_189_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_189,
        FIN => FIN_ANDGate_189,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_190 signals
    ANDGate_190: entity work.ANDGate_190
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_190
        output_190_Value => DecoderOutput_190_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_190,
        FIN => FIN_ANDGate_190,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_191 signals
    ANDGate_191: entity work.ANDGate_191
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderNOTInput_6
        m_input_NOT_6_Value => DecoderNOTInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_191
        output_191_Value => DecoderOutput_191_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_191,
        FIN => FIN_ANDGate_191,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_192 signals
    ANDGate_192: entity work.ANDGate_192
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_192
        output_192_Value => DecoderOutput_192_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_192,
        FIN => FIN_ANDGate_192,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_193 signals
    ANDGate_193: entity work.ANDGate_193
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_193
        output_193_Value => DecoderOutput_193_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_193,
        FIN => FIN_ANDGate_193,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_194 signals
    ANDGate_194: entity work.ANDGate_194
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_194
        output_194_Value => DecoderOutput_194_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_194,
        FIN => FIN_ANDGate_194,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_195 signals
    ANDGate_195: entity work.ANDGate_195
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_195
        output_195_Value => DecoderOutput_195_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_195,
        FIN => FIN_ANDGate_195,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_196 signals
    ANDGate_196: entity work.ANDGate_196
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_196
        output_196_Value => DecoderOutput_196_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_196,
        FIN => FIN_ANDGate_196,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_197 signals
    ANDGate_197: entity work.ANDGate_197
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_197
        output_197_Value => DecoderOutput_197_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_197,
        FIN => FIN_ANDGate_197,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_198 signals
    ANDGate_198: entity work.ANDGate_198
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_198
        output_198_Value => DecoderOutput_198_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_198,
        FIN => FIN_ANDGate_198,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_199 signals
    ANDGate_199: entity work.ANDGate_199
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_199
        output_199_Value => DecoderOutput_199_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_199,
        FIN => FIN_ANDGate_199,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_200 signals
    ANDGate_200: entity work.ANDGate_200
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_200
        output_200_Value => DecoderOutput_200_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_200,
        FIN => FIN_ANDGate_200,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_201 signals
    ANDGate_201: entity work.ANDGate_201
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_201
        output_201_Value => DecoderOutput_201_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_201,
        FIN => FIN_ANDGate_201,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_202 signals
    ANDGate_202: entity work.ANDGate_202
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_202
        output_202_Value => DecoderOutput_202_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_202,
        FIN => FIN_ANDGate_202,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_203 signals
    ANDGate_203: entity work.ANDGate_203
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_203
        output_203_Value => DecoderOutput_203_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_203,
        FIN => FIN_ANDGate_203,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_204 signals
    ANDGate_204: entity work.ANDGate_204
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_204
        output_204_Value => DecoderOutput_204_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_204,
        FIN => FIN_ANDGate_204,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_205 signals
    ANDGate_205: entity work.ANDGate_205
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_205
        output_205_Value => DecoderOutput_205_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_205,
        FIN => FIN_ANDGate_205,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_206 signals
    ANDGate_206: entity work.ANDGate_206
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_206
        output_206_Value => DecoderOutput_206_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_206,
        FIN => FIN_ANDGate_206,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_207 signals
    ANDGate_207: entity work.ANDGate_207
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_207
        output_207_Value => DecoderOutput_207_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_207,
        FIN => FIN_ANDGate_207,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_208 signals
    ANDGate_208: entity work.ANDGate_208
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_208
        output_208_Value => DecoderOutput_208_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_208,
        FIN => FIN_ANDGate_208,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_209 signals
    ANDGate_209: entity work.ANDGate_209
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_209
        output_209_Value => DecoderOutput_209_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_209,
        FIN => FIN_ANDGate_209,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_210 signals
    ANDGate_210: entity work.ANDGate_210
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_210
        output_210_Value => DecoderOutput_210_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_210,
        FIN => FIN_ANDGate_210,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_211 signals
    ANDGate_211: entity work.ANDGate_211
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_211
        output_211_Value => DecoderOutput_211_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_211,
        FIN => FIN_ANDGate_211,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_212 signals
    ANDGate_212: entity work.ANDGate_212
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_212
        output_212_Value => DecoderOutput_212_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_212,
        FIN => FIN_ANDGate_212,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_213 signals
    ANDGate_213: entity work.ANDGate_213
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_213
        output_213_Value => DecoderOutput_213_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_213,
        FIN => FIN_ANDGate_213,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_214 signals
    ANDGate_214: entity work.ANDGate_214
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_214
        output_214_Value => DecoderOutput_214_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_214,
        FIN => FIN_ANDGate_214,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_215 signals
    ANDGate_215: entity work.ANDGate_215
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_215
        output_215_Value => DecoderOutput_215_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_215,
        FIN => FIN_ANDGate_215,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_216 signals
    ANDGate_216: entity work.ANDGate_216
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_216
        output_216_Value => DecoderOutput_216_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_216,
        FIN => FIN_ANDGate_216,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_217 signals
    ANDGate_217: entity work.ANDGate_217
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_217
        output_217_Value => DecoderOutput_217_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_217,
        FIN => FIN_ANDGate_217,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_218 signals
    ANDGate_218: entity work.ANDGate_218
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_218
        output_218_Value => DecoderOutput_218_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_218,
        FIN => FIN_ANDGate_218,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_219 signals
    ANDGate_219: entity work.ANDGate_219
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_219
        output_219_Value => DecoderOutput_219_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_219,
        FIN => FIN_ANDGate_219,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_220 signals
    ANDGate_220: entity work.ANDGate_220
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_220
        output_220_Value => DecoderOutput_220_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_220,
        FIN => FIN_ANDGate_220,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_221 signals
    ANDGate_221: entity work.ANDGate_221
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_221
        output_221_Value => DecoderOutput_221_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_221,
        FIN => FIN_ANDGate_221,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_222 signals
    ANDGate_222: entity work.ANDGate_222
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_222
        output_222_Value => DecoderOutput_222_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_222,
        FIN => FIN_ANDGate_222,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_223 signals
    ANDGate_223: entity work.ANDGate_223
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderNOTInput_5
        m_input_NOT_5_Value => DecoderNOTInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_223
        output_223_Value => DecoderOutput_223_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_223,
        FIN => FIN_ANDGate_223,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_224 signals
    ANDGate_224: entity work.ANDGate_224
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_224
        output_224_Value => DecoderOutput_224_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_224,
        FIN => FIN_ANDGate_224,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_225 signals
    ANDGate_225: entity work.ANDGate_225
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_225
        output_225_Value => DecoderOutput_225_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_225,
        FIN => FIN_ANDGate_225,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_226 signals
    ANDGate_226: entity work.ANDGate_226
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_226
        output_226_Value => DecoderOutput_226_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_226,
        FIN => FIN_ANDGate_226,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_227 signals
    ANDGate_227: entity work.ANDGate_227
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_227
        output_227_Value => DecoderOutput_227_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_227,
        FIN => FIN_ANDGate_227,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_228 signals
    ANDGate_228: entity work.ANDGate_228
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_228
        output_228_Value => DecoderOutput_228_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_228,
        FIN => FIN_ANDGate_228,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_229 signals
    ANDGate_229: entity work.ANDGate_229
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_229
        output_229_Value => DecoderOutput_229_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_229,
        FIN => FIN_ANDGate_229,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_230 signals
    ANDGate_230: entity work.ANDGate_230
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_230
        output_230_Value => DecoderOutput_230_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_230,
        FIN => FIN_ANDGate_230,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_231 signals
    ANDGate_231: entity work.ANDGate_231
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_231
        output_231_Value => DecoderOutput_231_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_231,
        FIN => FIN_ANDGate_231,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_232 signals
    ANDGate_232: entity work.ANDGate_232
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_232
        output_232_Value => DecoderOutput_232_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_232,
        FIN => FIN_ANDGate_232,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_233 signals
    ANDGate_233: entity work.ANDGate_233
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_233
        output_233_Value => DecoderOutput_233_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_233,
        FIN => FIN_ANDGate_233,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_234 signals
    ANDGate_234: entity work.ANDGate_234
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_234
        output_234_Value => DecoderOutput_234_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_234,
        FIN => FIN_ANDGate_234,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_235 signals
    ANDGate_235: entity work.ANDGate_235
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_235
        output_235_Value => DecoderOutput_235_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_235,
        FIN => FIN_ANDGate_235,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_236 signals
    ANDGate_236: entity work.ANDGate_236
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_236
        output_236_Value => DecoderOutput_236_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_236,
        FIN => FIN_ANDGate_236,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_237 signals
    ANDGate_237: entity work.ANDGate_237
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_237
        output_237_Value => DecoderOutput_237_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_237,
        FIN => FIN_ANDGate_237,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_238 signals
    ANDGate_238: entity work.ANDGate_238
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_238
        output_238_Value => DecoderOutput_238_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_238,
        FIN => FIN_ANDGate_238,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_239 signals
    ANDGate_239: entity work.ANDGate_239
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderNOTInput_4
        m_input_NOT_4_Value => DecoderNOTInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_239
        output_239_Value => DecoderOutput_239_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_239,
        FIN => FIN_ANDGate_239,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_240 signals
    ANDGate_240: entity work.ANDGate_240
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_240
        output_240_Value => DecoderOutput_240_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_240,
        FIN => FIN_ANDGate_240,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_241 signals
    ANDGate_241: entity work.ANDGate_241
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_241
        output_241_Value => DecoderOutput_241_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_241,
        FIN => FIN_ANDGate_241,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_242 signals
    ANDGate_242: entity work.ANDGate_242
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_242
        output_242_Value => DecoderOutput_242_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_242,
        FIN => FIN_ANDGate_242,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_243 signals
    ANDGate_243: entity work.ANDGate_243
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_243
        output_243_Value => DecoderOutput_243_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_243,
        FIN => FIN_ANDGate_243,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_244 signals
    ANDGate_244: entity work.ANDGate_244
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_244
        output_244_Value => DecoderOutput_244_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_244,
        FIN => FIN_ANDGate_244,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_245 signals
    ANDGate_245: entity work.ANDGate_245
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_245
        output_245_Value => DecoderOutput_245_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_245,
        FIN => FIN_ANDGate_245,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_246 signals
    ANDGate_246: entity work.ANDGate_246
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_246
        output_246_Value => DecoderOutput_246_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_246,
        FIN => FIN_ANDGate_246,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_247 signals
    ANDGate_247: entity work.ANDGate_247
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderNOTInput_3
        m_input_NOT_3_Value => DecoderNOTInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_247
        output_247_Value => DecoderOutput_247_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_247,
        FIN => FIN_ANDGate_247,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_248 signals
    ANDGate_248: entity work.ANDGate_248
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_248
        output_248_Value => DecoderOutput_248_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_248,
        FIN => FIN_ANDGate_248,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_249 signals
    ANDGate_249: entity work.ANDGate_249
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_249
        output_249_Value => DecoderOutput_249_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_249,
        FIN => FIN_ANDGate_249,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_250 signals
    ANDGate_250: entity work.ANDGate_250
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_250
        output_250_Value => DecoderOutput_250_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_250,
        FIN => FIN_ANDGate_250,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_251 signals
    ANDGate_251: entity work.ANDGate_251
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderNOTInput_2
        m_input_NOT_2_Value => DecoderNOTInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_251
        output_251_Value => DecoderOutput_251_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_251,
        FIN => FIN_ANDGate_251,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_252 signals
    ANDGate_252: entity work.ANDGate_252
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_252
        output_252_Value => DecoderOutput_252_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_252,
        FIN => FIN_ANDGate_252,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_253 signals
    ANDGate_253: entity work.ANDGate_253
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderNOTInput_1
        m_input_NOT_1_Value => DecoderNOTInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_253
        output_253_Value => DecoderOutput_253_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_253,
        FIN => FIN_ANDGate_253,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_254 signals
    ANDGate_254: entity work.ANDGate_254
    port map (
        -- Input bus DecoderNOTInput_0
        m_input_NOT_0_Value => DecoderNOTInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_254
        output_254_Value => DecoderOutput_254_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_254,
        FIN => FIN_ANDGate_254,
        ENB => ENB,
        RST => RST
    );


    -- Entity  ANDGate_255 signals
    ANDGate_255: entity work.ANDGate_255
    port map (
        -- Input bus DecoderInput_0
        m_input_0_Value => DecoderInput_0_Value,


        -- Input bus DecoderInput_1
        m_input_1_Value => DecoderInput_1_Value,


        -- Input bus DecoderInput_2
        m_input_2_Value => DecoderInput_2_Value,


        -- Input bus DecoderInput_3
        m_input_3_Value => DecoderInput_3_Value,


        -- Input bus DecoderInput_4
        m_input_4_Value => DecoderInput_4_Value,


        -- Input bus DecoderInput_5
        m_input_5_Value => DecoderInput_5_Value,


        -- Input bus DecoderInput_6
        m_input_6_Value => DecoderInput_6_Value,


        -- Input bus DecoderInput_7
        m_input_7_Value => DecoderInput_7_Value,


        -- Output bus DecoderOutput_255
        output_255_Value => DecoderOutput_255_Value,



        CLK => CLK,
        RDY => RDY_ANDGate_255,
        FIN => FIN_ANDGate_255,
        ENB => ENB,
        RST => RST
    );


    -- Connect ready signals
    RDY_NOTGate_0 <= RDY;
    RDY_NOTGate_1 <= RDY;
    RDY_NOTGate_2 <= RDY;
    RDY_NOTGate_3 <= RDY;
    RDY_NOTGate_4 <= RDY;
    RDY_NOTGate_5 <= RDY;
    RDY_NOTGate_6 <= RDY;
    RDY_NOTGate_7 <= RDY;
    -- Setup the RDY signal for ANDGate_0
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_0 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_1
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_1 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_2
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_2 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_3
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_6 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_3 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_4
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_4 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_5
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_5 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_6
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_6 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_7
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_4 AND FIN_NOTGate_3 = FIN_NOTGate_5 AND FIN_NOTGate_3 = FIN_NOTGate_6 AND FIN_NOTGate_3 = FIN_NOTGate_7 then
        RDY_ANDGate_7 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_8
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_8 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_9
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_9 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_10
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_10 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_11
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_6 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_11 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_12
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_12 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_13
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_13 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_14
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_14 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_15
    process(
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_4 = FIN_NOTGate_5 AND FIN_NOTGate_4 = FIN_NOTGate_6 AND FIN_NOTGate_4 = FIN_NOTGate_7 then
        RDY_ANDGate_15 <= FIN_NOTGate_4;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_16
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_16 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_17
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_17 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_18
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_18 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_19
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_6 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_19 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_20
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_20 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_21
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_21 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_22
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_22 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_23
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_5 AND FIN_NOTGate_3 = FIN_NOTGate_6 AND FIN_NOTGate_3 = FIN_NOTGate_7 then
        RDY_ANDGate_23 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_24
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_24 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_25
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_25 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_26
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_26 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_27
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_6 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_27 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_28
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_28 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_29
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_29 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_30
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_30 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_31
    process(
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_5 = FIN_NOTGate_6 AND FIN_NOTGate_5 = FIN_NOTGate_7 then
        RDY_ANDGate_31 <= FIN_NOTGate_5;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_32
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_32 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_33
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_33 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_34
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_34 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_35
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_6 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_35 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_36
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_36 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_37
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_37 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_38
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_38 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_39
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_4 AND FIN_NOTGate_3 = FIN_NOTGate_6 AND FIN_NOTGate_3 = FIN_NOTGate_7 then
        RDY_ANDGate_39 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_40
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_40 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_41
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_41 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_42
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_42 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_43
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_6 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_43 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_44
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_44 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_45
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_45 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_46
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_46 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_47
    process(
      FIN_NOTGate_4, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_4 = FIN_NOTGate_6 AND FIN_NOTGate_4 = FIN_NOTGate_7 then
        RDY_ANDGate_47 <= FIN_NOTGate_4;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_48
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_48 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_49
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_49 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_50
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_50 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_51
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_6 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_51 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_52
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_52 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_53
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_53 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_54
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_54 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_55
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_6 AND FIN_NOTGate_3 = FIN_NOTGate_7 then
        RDY_ANDGate_55 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_56
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_56 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_57
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_57 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_58
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_58 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_59
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_6 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_59 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_60
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_60 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_61
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_6 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_61 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_62
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_62 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_63
    process(
      FIN_NOTGate_6, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_6 = FIN_NOTGate_7 then
        RDY_ANDGate_63 <= FIN_NOTGate_6;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_64
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_64 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_65
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_65 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_66
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_66 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_67
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_67 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_68
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_68 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_69
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_69 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_70
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_70 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_71
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_4 AND FIN_NOTGate_3 = FIN_NOTGate_5 AND FIN_NOTGate_3 = FIN_NOTGate_7 then
        RDY_ANDGate_71 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_72
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_72 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_73
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_73 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_74
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_74 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_75
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_75 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_76
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_76 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_77
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_77 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_78
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_78 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_79
    process(
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_4 = FIN_NOTGate_5 AND FIN_NOTGate_4 = FIN_NOTGate_7 then
        RDY_ANDGate_79 <= FIN_NOTGate_4;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_80
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_80 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_81
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_81 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_82
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_82 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_83
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_83 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_84
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_84 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_85
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_85 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_86
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_86 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_87
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_5 AND FIN_NOTGate_3 = FIN_NOTGate_7 then
        RDY_ANDGate_87 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_88
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_88 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_89
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_89 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_90
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_90 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_91
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_91 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_92
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_92 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_93
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_93 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_94
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_94 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_95
    process(
      FIN_NOTGate_5, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_5 = FIN_NOTGate_7 then
        RDY_ANDGate_95 <= FIN_NOTGate_5;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_96
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_96 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_97
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_97 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_98
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_98 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_99
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_99 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_100
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_100 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_101
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_101 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_102
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_102 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_103
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_4 AND FIN_NOTGate_3 = FIN_NOTGate_7 then
        RDY_ANDGate_103 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_104
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_104 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_105
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_105 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_106
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_106 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_107
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_107 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_108
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_108 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_109
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_109 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_110
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_110 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_111
    process(
      FIN_NOTGate_4, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_4 = FIN_NOTGate_7 then
        RDY_ANDGate_111 <= FIN_NOTGate_4;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_112
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_112 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_113
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_113 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_114
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_114 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_115
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_115 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_116
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_116 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_117
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_117 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_118
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_118 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_119
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_7 then
        RDY_ANDGate_119 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_120
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_120 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_121
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_121 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_122
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_122 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_123
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_7 then
        RDY_ANDGate_123 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_124
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_124 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_125
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_7 then
        RDY_ANDGate_125 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_126
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_7
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_7 then
        RDY_ANDGate_126 <= FIN_NOTGate_0;
      end if;
    end process;
    RDY_ANDGate_127 <= FIN_NOTGate_7;
    -- Setup the RDY signal for ANDGate_128
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_128 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_129
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_129 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_130
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_130 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_131
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_6 then
        RDY_ANDGate_131 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_132
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_132 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_133
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_133 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_134
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_134 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_135
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_4 AND FIN_NOTGate_3 = FIN_NOTGate_5 AND FIN_NOTGate_3 = FIN_NOTGate_6 then
        RDY_ANDGate_135 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_136
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_136 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_137
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_137 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_138
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_138 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_139
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_6 then
        RDY_ANDGate_139 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_140
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_140 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_141
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_141 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_142
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_142 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_143
    process(
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_4 = FIN_NOTGate_5 AND FIN_NOTGate_4 = FIN_NOTGate_6 then
        RDY_ANDGate_143 <= FIN_NOTGate_4;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_144
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_144 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_145
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_145 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_146
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_146 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_147
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_6 then
        RDY_ANDGate_147 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_148
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_148 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_149
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_149 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_150
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_150 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_151
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_5 AND FIN_NOTGate_3 = FIN_NOTGate_6 then
        RDY_ANDGate_151 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_152
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_152 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_153
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_153 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_154
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_154 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_155
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_5 AND FIN_NOTGate_2 = FIN_NOTGate_6 then
        RDY_ANDGate_155 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_156
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_156 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_157
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_5 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_157 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_158
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_158 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_159
    process(
      FIN_NOTGate_5, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_5 = FIN_NOTGate_6 then
        RDY_ANDGate_159 <= FIN_NOTGate_5;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_160
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_160 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_161
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_161 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_162
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_162 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_163
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_6 then
        RDY_ANDGate_163 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_164
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_164 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_165
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_165 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_166
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_166 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_167
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_4 AND FIN_NOTGate_3 = FIN_NOTGate_6 then
        RDY_ANDGate_167 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_168
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_168 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_169
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_169 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_170
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_170 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_171
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_6 then
        RDY_ANDGate_171 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_172
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_172 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_173
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_173 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_174
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_174 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_175
    process(
      FIN_NOTGate_4, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_4 = FIN_NOTGate_6 then
        RDY_ANDGate_175 <= FIN_NOTGate_4;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_176
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_176 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_177
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_177 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_178
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_178 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_179
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_6 then
        RDY_ANDGate_179 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_180
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_180 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_181
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_181 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_182
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_182 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_183
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_6 then
        RDY_ANDGate_183 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_184
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_184 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_185
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_185 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_186
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_186 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_187
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_6 then
        RDY_ANDGate_187 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_188
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_188 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_189
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_6 then
        RDY_ANDGate_189 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_190
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_6
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_6 then
        RDY_ANDGate_190 <= FIN_NOTGate_0;
      end if;
    end process;
    RDY_ANDGate_191 <= FIN_NOTGate_6;
    -- Setup the RDY signal for ANDGate_192
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_192 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_193
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 then
        RDY_ANDGate_193 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_194
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_194 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_195
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_5 then
        RDY_ANDGate_195 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_196
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_196 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_197
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 then
        RDY_ANDGate_197 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_198
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_198 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_199
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_4 AND FIN_NOTGate_3 = FIN_NOTGate_5 then
        RDY_ANDGate_199 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_200
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_200 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_201
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 then
        RDY_ANDGate_201 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_202
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_202 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_203
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_4 AND FIN_NOTGate_2 = FIN_NOTGate_5 then
        RDY_ANDGate_203 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_204
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_204 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_205
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_4 AND FIN_NOTGate_1 = FIN_NOTGate_5 then
        RDY_ANDGate_205 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_206
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_206 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_207
    process(
      FIN_NOTGate_4, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_4 = FIN_NOTGate_5 then
        RDY_ANDGate_207 <= FIN_NOTGate_4;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_208
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_208 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_209
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_5 then
        RDY_ANDGate_209 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_210
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_210 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_211
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_5 then
        RDY_ANDGate_211 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_212
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_212 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_213
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_5 then
        RDY_ANDGate_213 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_214
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_214 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_215
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_5 then
        RDY_ANDGate_215 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_216
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_216 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_217
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_5 then
        RDY_ANDGate_217 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_218
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_218 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_219
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_5 then
        RDY_ANDGate_219 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_220
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_220 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_221
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_5 then
        RDY_ANDGate_221 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_222
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_5
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_5 then
        RDY_ANDGate_222 <= FIN_NOTGate_0;
      end if;
    end process;
    RDY_ANDGate_223 <= FIN_NOTGate_5;
    -- Setup the RDY signal for ANDGate_224
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 then
        RDY_ANDGate_224 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_225
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 then
        RDY_ANDGate_225 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_226
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 then
        RDY_ANDGate_226 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_227
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 AND FIN_NOTGate_2 = FIN_NOTGate_4 then
        RDY_ANDGate_227 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_228
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 then
        RDY_ANDGate_228 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_229
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 AND FIN_NOTGate_1 = FIN_NOTGate_4 then
        RDY_ANDGate_229 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_230
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 then
        RDY_ANDGate_230 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_231
    process(
      FIN_NOTGate_3, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_3 = FIN_NOTGate_4 then
        RDY_ANDGate_231 <= FIN_NOTGate_3;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_232
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 then
        RDY_ANDGate_232 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_233
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_4 then
        RDY_ANDGate_233 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_234
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_4 then
        RDY_ANDGate_234 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_235
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_4 then
        RDY_ANDGate_235 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_236
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_4 then
        RDY_ANDGate_236 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_237
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_4 then
        RDY_ANDGate_237 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_238
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_4
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_4 then
        RDY_ANDGate_238 <= FIN_NOTGate_0;
      end if;
    end process;
    RDY_ANDGate_239 <= FIN_NOTGate_4;
    -- Setup the RDY signal for ANDGate_240
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 then
        RDY_ANDGate_240 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_241
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 AND FIN_NOTGate_1 = FIN_NOTGate_3 then
        RDY_ANDGate_241 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_242
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 then
        RDY_ANDGate_242 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_243
    process(
      FIN_NOTGate_2, 
      FIN_NOTGate_3
    )
    begin
      if FIN_NOTGate_2 = FIN_NOTGate_3 then
        RDY_ANDGate_243 <= FIN_NOTGate_2;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_244
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_3
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_3 then
        RDY_ANDGate_244 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_245
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_3
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_3 then
        RDY_ANDGate_245 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_246
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_3
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_3 then
        RDY_ANDGate_246 <= FIN_NOTGate_0;
      end if;
    end process;
    RDY_ANDGate_247 <= FIN_NOTGate_3;
    -- Setup the RDY signal for ANDGate_248
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 then
        RDY_ANDGate_248 <= FIN_NOTGate_0;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_249
    process(
      FIN_NOTGate_1, 
      FIN_NOTGate_2
    )
    begin
      if FIN_NOTGate_1 = FIN_NOTGate_2 then
        RDY_ANDGate_249 <= FIN_NOTGate_1;
      end if;
    end process;
    -- Setup the RDY signal for ANDGate_250
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_2
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_2 then
        RDY_ANDGate_250 <= FIN_NOTGate_0;
      end if;
    end process;
    RDY_ANDGate_251 <= FIN_NOTGate_2;
    -- Setup the RDY signal for ANDGate_252
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 then
        RDY_ANDGate_252 <= FIN_NOTGate_0;
      end if;
    end process;
    RDY_ANDGate_253 <= FIN_NOTGate_1;
    RDY_ANDGate_254 <= FIN_NOTGate_0;
    RDY_ANDGate_255 <= RDY;

    -- Setup the FIN feedback signals
    process(
      FIN_NOTGate_0, 
      FIN_NOTGate_1, 
      FIN_NOTGate_2, 
      FIN_NOTGate_3, 
      FIN_NOTGate_4, 
      FIN_NOTGate_5, 
      FIN_NOTGate_6, 
      FIN_NOTGate_7, 
      FIN_ANDGate_0, 
      FIN_ANDGate_1, 
      FIN_ANDGate_2, 
      FIN_ANDGate_3, 
      FIN_ANDGate_4, 
      FIN_ANDGate_5, 
      FIN_ANDGate_6, 
      FIN_ANDGate_7, 
      FIN_ANDGate_8, 
      FIN_ANDGate_9, 
      FIN_ANDGate_10, 
      FIN_ANDGate_11, 
      FIN_ANDGate_12, 
      FIN_ANDGate_13, 
      FIN_ANDGate_14, 
      FIN_ANDGate_15, 
      FIN_ANDGate_16, 
      FIN_ANDGate_17, 
      FIN_ANDGate_18, 
      FIN_ANDGate_19, 
      FIN_ANDGate_20, 
      FIN_ANDGate_21, 
      FIN_ANDGate_22, 
      FIN_ANDGate_23, 
      FIN_ANDGate_24, 
      FIN_ANDGate_25, 
      FIN_ANDGate_26, 
      FIN_ANDGate_27, 
      FIN_ANDGate_28, 
      FIN_ANDGate_29, 
      FIN_ANDGate_30, 
      FIN_ANDGate_31, 
      FIN_ANDGate_32, 
      FIN_ANDGate_33, 
      FIN_ANDGate_34, 
      FIN_ANDGate_35, 
      FIN_ANDGate_36, 
      FIN_ANDGate_37, 
      FIN_ANDGate_38, 
      FIN_ANDGate_39, 
      FIN_ANDGate_40, 
      FIN_ANDGate_41, 
      FIN_ANDGate_42, 
      FIN_ANDGate_43, 
      FIN_ANDGate_44, 
      FIN_ANDGate_45, 
      FIN_ANDGate_46, 
      FIN_ANDGate_47, 
      FIN_ANDGate_48, 
      FIN_ANDGate_49, 
      FIN_ANDGate_50, 
      FIN_ANDGate_51, 
      FIN_ANDGate_52, 
      FIN_ANDGate_53, 
      FIN_ANDGate_54, 
      FIN_ANDGate_55, 
      FIN_ANDGate_56, 
      FIN_ANDGate_57, 
      FIN_ANDGate_58, 
      FIN_ANDGate_59, 
      FIN_ANDGate_60, 
      FIN_ANDGate_61, 
      FIN_ANDGate_62, 
      FIN_ANDGate_63, 
      FIN_ANDGate_64, 
      FIN_ANDGate_65, 
      FIN_ANDGate_66, 
      FIN_ANDGate_67, 
      FIN_ANDGate_68, 
      FIN_ANDGate_69, 
      FIN_ANDGate_70, 
      FIN_ANDGate_71, 
      FIN_ANDGate_72, 
      FIN_ANDGate_73, 
      FIN_ANDGate_74, 
      FIN_ANDGate_75, 
      FIN_ANDGate_76, 
      FIN_ANDGate_77, 
      FIN_ANDGate_78, 
      FIN_ANDGate_79, 
      FIN_ANDGate_80, 
      FIN_ANDGate_81, 
      FIN_ANDGate_82, 
      FIN_ANDGate_83, 
      FIN_ANDGate_84, 
      FIN_ANDGate_85, 
      FIN_ANDGate_86, 
      FIN_ANDGate_87, 
      FIN_ANDGate_88, 
      FIN_ANDGate_89, 
      FIN_ANDGate_90, 
      FIN_ANDGate_91, 
      FIN_ANDGate_92, 
      FIN_ANDGate_93, 
      FIN_ANDGate_94, 
      FIN_ANDGate_95, 
      FIN_ANDGate_96, 
      FIN_ANDGate_97, 
      FIN_ANDGate_98, 
      FIN_ANDGate_99, 
      FIN_ANDGate_100, 
      FIN_ANDGate_101, 
      FIN_ANDGate_102, 
      FIN_ANDGate_103, 
      FIN_ANDGate_104, 
      FIN_ANDGate_105, 
      FIN_ANDGate_106, 
      FIN_ANDGate_107, 
      FIN_ANDGate_108, 
      FIN_ANDGate_109, 
      FIN_ANDGate_110, 
      FIN_ANDGate_111, 
      FIN_ANDGate_112, 
      FIN_ANDGate_113, 
      FIN_ANDGate_114, 
      FIN_ANDGate_115, 
      FIN_ANDGate_116, 
      FIN_ANDGate_117, 
      FIN_ANDGate_118, 
      FIN_ANDGate_119, 
      FIN_ANDGate_120, 
      FIN_ANDGate_121, 
      FIN_ANDGate_122, 
      FIN_ANDGate_123, 
      FIN_ANDGate_124, 
      FIN_ANDGate_125, 
      FIN_ANDGate_126, 
      FIN_ANDGate_127, 
      FIN_ANDGate_128, 
      FIN_ANDGate_129, 
      FIN_ANDGate_130, 
      FIN_ANDGate_131, 
      FIN_ANDGate_132, 
      FIN_ANDGate_133, 
      FIN_ANDGate_134, 
      FIN_ANDGate_135, 
      FIN_ANDGate_136, 
      FIN_ANDGate_137, 
      FIN_ANDGate_138, 
      FIN_ANDGate_139, 
      FIN_ANDGate_140, 
      FIN_ANDGate_141, 
      FIN_ANDGate_142, 
      FIN_ANDGate_143, 
      FIN_ANDGate_144, 
      FIN_ANDGate_145, 
      FIN_ANDGate_146, 
      FIN_ANDGate_147, 
      FIN_ANDGate_148, 
      FIN_ANDGate_149, 
      FIN_ANDGate_150, 
      FIN_ANDGate_151, 
      FIN_ANDGate_152, 
      FIN_ANDGate_153, 
      FIN_ANDGate_154, 
      FIN_ANDGate_155, 
      FIN_ANDGate_156, 
      FIN_ANDGate_157, 
      FIN_ANDGate_158, 
      FIN_ANDGate_159, 
      FIN_ANDGate_160, 
      FIN_ANDGate_161, 
      FIN_ANDGate_162, 
      FIN_ANDGate_163, 
      FIN_ANDGate_164, 
      FIN_ANDGate_165, 
      FIN_ANDGate_166, 
      FIN_ANDGate_167, 
      FIN_ANDGate_168, 
      FIN_ANDGate_169, 
      FIN_ANDGate_170, 
      FIN_ANDGate_171, 
      FIN_ANDGate_172, 
      FIN_ANDGate_173, 
      FIN_ANDGate_174, 
      FIN_ANDGate_175, 
      FIN_ANDGate_176, 
      FIN_ANDGate_177, 
      FIN_ANDGate_178, 
      FIN_ANDGate_179, 
      FIN_ANDGate_180, 
      FIN_ANDGate_181, 
      FIN_ANDGate_182, 
      FIN_ANDGate_183, 
      FIN_ANDGate_184, 
      FIN_ANDGate_185, 
      FIN_ANDGate_186, 
      FIN_ANDGate_187, 
      FIN_ANDGate_188, 
      FIN_ANDGate_189, 
      FIN_ANDGate_190, 
      FIN_ANDGate_191, 
      FIN_ANDGate_192, 
      FIN_ANDGate_193, 
      FIN_ANDGate_194, 
      FIN_ANDGate_195, 
      FIN_ANDGate_196, 
      FIN_ANDGate_197, 
      FIN_ANDGate_198, 
      FIN_ANDGate_199, 
      FIN_ANDGate_200, 
      FIN_ANDGate_201, 
      FIN_ANDGate_202, 
      FIN_ANDGate_203, 
      FIN_ANDGate_204, 
      FIN_ANDGate_205, 
      FIN_ANDGate_206, 
      FIN_ANDGate_207, 
      FIN_ANDGate_208, 
      FIN_ANDGate_209, 
      FIN_ANDGate_210, 
      FIN_ANDGate_211, 
      FIN_ANDGate_212, 
      FIN_ANDGate_213, 
      FIN_ANDGate_214, 
      FIN_ANDGate_215, 
      FIN_ANDGate_216, 
      FIN_ANDGate_217, 
      FIN_ANDGate_218, 
      FIN_ANDGate_219, 
      FIN_ANDGate_220, 
      FIN_ANDGate_221, 
      FIN_ANDGate_222, 
      FIN_ANDGate_223, 
      FIN_ANDGate_224, 
      FIN_ANDGate_225, 
      FIN_ANDGate_226, 
      FIN_ANDGate_227, 
      FIN_ANDGate_228, 
      FIN_ANDGate_229, 
      FIN_ANDGate_230, 
      FIN_ANDGate_231, 
      FIN_ANDGate_232, 
      FIN_ANDGate_233, 
      FIN_ANDGate_234, 
      FIN_ANDGate_235, 
      FIN_ANDGate_236, 
      FIN_ANDGate_237, 
      FIN_ANDGate_238, 
      FIN_ANDGate_239, 
      FIN_ANDGate_240, 
      FIN_ANDGate_241, 
      FIN_ANDGate_242, 
      FIN_ANDGate_243, 
      FIN_ANDGate_244, 
      FIN_ANDGate_245, 
      FIN_ANDGate_246, 
      FIN_ANDGate_247, 
      FIN_ANDGate_248, 
      FIN_ANDGate_249, 
      FIN_ANDGate_250, 
      FIN_ANDGate_251, 
      FIN_ANDGate_252, 
      FIN_ANDGate_253, 
      FIN_ANDGate_254, 
      FIN_ANDGate_255
    )
    begin
      if FIN_NOTGate_0 = FIN_NOTGate_1 AND FIN_NOTGate_0 = FIN_NOTGate_2 AND FIN_NOTGate_0 = FIN_NOTGate_3 AND FIN_NOTGate_0 = FIN_NOTGate_4 AND FIN_NOTGate_0 = FIN_NOTGate_5 AND FIN_NOTGate_0 = FIN_NOTGate_6 AND FIN_NOTGate_0 = FIN_NOTGate_7 AND FIN_NOTGate_0 = FIN_ANDGate_0 AND FIN_NOTGate_0 = FIN_ANDGate_1 AND FIN_NOTGate_0 = FIN_ANDGate_2 AND FIN_NOTGate_0 = FIN_ANDGate_3 AND FIN_NOTGate_0 = FIN_ANDGate_4 AND FIN_NOTGate_0 = FIN_ANDGate_5 AND FIN_NOTGate_0 = FIN_ANDGate_6 AND FIN_NOTGate_0 = FIN_ANDGate_7 AND FIN_NOTGate_0 = FIN_ANDGate_8 AND FIN_NOTGate_0 = FIN_ANDGate_9 AND FIN_NOTGate_0 = FIN_ANDGate_10 AND FIN_NOTGate_0 = FIN_ANDGate_11 AND FIN_NOTGate_0 = FIN_ANDGate_12 AND FIN_NOTGate_0 = FIN_ANDGate_13 AND FIN_NOTGate_0 = FIN_ANDGate_14 AND FIN_NOTGate_0 = FIN_ANDGate_15 AND FIN_NOTGate_0 = FIN_ANDGate_16 AND FIN_NOTGate_0 = FIN_ANDGate_17 AND FIN_NOTGate_0 = FIN_ANDGate_18 AND FIN_NOTGate_0 = FIN_ANDGate_19 AND FIN_NOTGate_0 = FIN_ANDGate_20 AND FIN_NOTGate_0 = FIN_ANDGate_21 AND FIN_NOTGate_0 = FIN_ANDGate_22 AND FIN_NOTGate_0 = FIN_ANDGate_23 AND FIN_NOTGate_0 = FIN_ANDGate_24 AND FIN_NOTGate_0 = FIN_ANDGate_25 AND FIN_NOTGate_0 = FIN_ANDGate_26 AND FIN_NOTGate_0 = FIN_ANDGate_27 AND FIN_NOTGate_0 = FIN_ANDGate_28 AND FIN_NOTGate_0 = FIN_ANDGate_29 AND FIN_NOTGate_0 = FIN_ANDGate_30 AND FIN_NOTGate_0 = FIN_ANDGate_31 AND FIN_NOTGate_0 = FIN_ANDGate_32 AND FIN_NOTGate_0 = FIN_ANDGate_33 AND FIN_NOTGate_0 = FIN_ANDGate_34 AND FIN_NOTGate_0 = FIN_ANDGate_35 AND FIN_NOTGate_0 = FIN_ANDGate_36 AND FIN_NOTGate_0 = FIN_ANDGate_37 AND FIN_NOTGate_0 = FIN_ANDGate_38 AND FIN_NOTGate_0 = FIN_ANDGate_39 AND FIN_NOTGate_0 = FIN_ANDGate_40 AND FIN_NOTGate_0 = FIN_ANDGate_41 AND FIN_NOTGate_0 = FIN_ANDGate_42 AND FIN_NOTGate_0 = FIN_ANDGate_43 AND FIN_NOTGate_0 = FIN_ANDGate_44 AND FIN_NOTGate_0 = FIN_ANDGate_45 AND FIN_NOTGate_0 = FIN_ANDGate_46 AND FIN_NOTGate_0 = FIN_ANDGate_47 AND FIN_NOTGate_0 = FIN_ANDGate_48 AND FIN_NOTGate_0 = FIN_ANDGate_49 AND FIN_NOTGate_0 = FIN_ANDGate_50 AND FIN_NOTGate_0 = FIN_ANDGate_51 AND FIN_NOTGate_0 = FIN_ANDGate_52 AND FIN_NOTGate_0 = FIN_ANDGate_53 AND FIN_NOTGate_0 = FIN_ANDGate_54 AND FIN_NOTGate_0 = FIN_ANDGate_55 AND FIN_NOTGate_0 = FIN_ANDGate_56 AND FIN_NOTGate_0 = FIN_ANDGate_57 AND FIN_NOTGate_0 = FIN_ANDGate_58 AND FIN_NOTGate_0 = FIN_ANDGate_59 AND FIN_NOTGate_0 = FIN_ANDGate_60 AND FIN_NOTGate_0 = FIN_ANDGate_61 AND FIN_NOTGate_0 = FIN_ANDGate_62 AND FIN_NOTGate_0 = FIN_ANDGate_63 AND FIN_NOTGate_0 = FIN_ANDGate_64 AND FIN_NOTGate_0 = FIN_ANDGate_65 AND FIN_NOTGate_0 = FIN_ANDGate_66 AND FIN_NOTGate_0 = FIN_ANDGate_67 AND FIN_NOTGate_0 = FIN_ANDGate_68 AND FIN_NOTGate_0 = FIN_ANDGate_69 AND FIN_NOTGate_0 = FIN_ANDGate_70 AND FIN_NOTGate_0 = FIN_ANDGate_71 AND FIN_NOTGate_0 = FIN_ANDGate_72 AND FIN_NOTGate_0 = FIN_ANDGate_73 AND FIN_NOTGate_0 = FIN_ANDGate_74 AND FIN_NOTGate_0 = FIN_ANDGate_75 AND FIN_NOTGate_0 = FIN_ANDGate_76 AND FIN_NOTGate_0 = FIN_ANDGate_77 AND FIN_NOTGate_0 = FIN_ANDGate_78 AND FIN_NOTGate_0 = FIN_ANDGate_79 AND FIN_NOTGate_0 = FIN_ANDGate_80 AND FIN_NOTGate_0 = FIN_ANDGate_81 AND FIN_NOTGate_0 = FIN_ANDGate_82 AND FIN_NOTGate_0 = FIN_ANDGate_83 AND FIN_NOTGate_0 = FIN_ANDGate_84 AND FIN_NOTGate_0 = FIN_ANDGate_85 AND FIN_NOTGate_0 = FIN_ANDGate_86 AND FIN_NOTGate_0 = FIN_ANDGate_87 AND FIN_NOTGate_0 = FIN_ANDGate_88 AND FIN_NOTGate_0 = FIN_ANDGate_89 AND FIN_NOTGate_0 = FIN_ANDGate_90 AND FIN_NOTGate_0 = FIN_ANDGate_91 AND FIN_NOTGate_0 = FIN_ANDGate_92 AND FIN_NOTGate_0 = FIN_ANDGate_93 AND FIN_NOTGate_0 = FIN_ANDGate_94 AND FIN_NOTGate_0 = FIN_ANDGate_95 AND FIN_NOTGate_0 = FIN_ANDGate_96 AND FIN_NOTGate_0 = FIN_ANDGate_97 AND FIN_NOTGate_0 = FIN_ANDGate_98 AND FIN_NOTGate_0 = FIN_ANDGate_99 AND FIN_NOTGate_0 = FIN_ANDGate_100 AND FIN_NOTGate_0 = FIN_ANDGate_101 AND FIN_NOTGate_0 = FIN_ANDGate_102 AND FIN_NOTGate_0 = FIN_ANDGate_103 AND FIN_NOTGate_0 = FIN_ANDGate_104 AND FIN_NOTGate_0 = FIN_ANDGate_105 AND FIN_NOTGate_0 = FIN_ANDGate_106 AND FIN_NOTGate_0 = FIN_ANDGate_107 AND FIN_NOTGate_0 = FIN_ANDGate_108 AND FIN_NOTGate_0 = FIN_ANDGate_109 AND FIN_NOTGate_0 = FIN_ANDGate_110 AND FIN_NOTGate_0 = FIN_ANDGate_111 AND FIN_NOTGate_0 = FIN_ANDGate_112 AND FIN_NOTGate_0 = FIN_ANDGate_113 AND FIN_NOTGate_0 = FIN_ANDGate_114 AND FIN_NOTGate_0 = FIN_ANDGate_115 AND FIN_NOTGate_0 = FIN_ANDGate_116 AND FIN_NOTGate_0 = FIN_ANDGate_117 AND FIN_NOTGate_0 = FIN_ANDGate_118 AND FIN_NOTGate_0 = FIN_ANDGate_119 AND FIN_NOTGate_0 = FIN_ANDGate_120 AND FIN_NOTGate_0 = FIN_ANDGate_121 AND FIN_NOTGate_0 = FIN_ANDGate_122 AND FIN_NOTGate_0 = FIN_ANDGate_123 AND FIN_NOTGate_0 = FIN_ANDGate_124 AND FIN_NOTGate_0 = FIN_ANDGate_125 AND FIN_NOTGate_0 = FIN_ANDGate_126 AND FIN_NOTGate_0 = FIN_ANDGate_127 AND FIN_NOTGate_0 = FIN_ANDGate_128 AND FIN_NOTGate_0 = FIN_ANDGate_129 AND FIN_NOTGate_0 = FIN_ANDGate_130 AND FIN_NOTGate_0 = FIN_ANDGate_131 AND FIN_NOTGate_0 = FIN_ANDGate_132 AND FIN_NOTGate_0 = FIN_ANDGate_133 AND FIN_NOTGate_0 = FIN_ANDGate_134 AND FIN_NOTGate_0 = FIN_ANDGate_135 AND FIN_NOTGate_0 = FIN_ANDGate_136 AND FIN_NOTGate_0 = FIN_ANDGate_137 AND FIN_NOTGate_0 = FIN_ANDGate_138 AND FIN_NOTGate_0 = FIN_ANDGate_139 AND FIN_NOTGate_0 = FIN_ANDGate_140 AND FIN_NOTGate_0 = FIN_ANDGate_141 AND FIN_NOTGate_0 = FIN_ANDGate_142 AND FIN_NOTGate_0 = FIN_ANDGate_143 AND FIN_NOTGate_0 = FIN_ANDGate_144 AND FIN_NOTGate_0 = FIN_ANDGate_145 AND FIN_NOTGate_0 = FIN_ANDGate_146 AND FIN_NOTGate_0 = FIN_ANDGate_147 AND FIN_NOTGate_0 = FIN_ANDGate_148 AND FIN_NOTGate_0 = FIN_ANDGate_149 AND FIN_NOTGate_0 = FIN_ANDGate_150 AND FIN_NOTGate_0 = FIN_ANDGate_151 AND FIN_NOTGate_0 = FIN_ANDGate_152 AND FIN_NOTGate_0 = FIN_ANDGate_153 AND FIN_NOTGate_0 = FIN_ANDGate_154 AND FIN_NOTGate_0 = FIN_ANDGate_155 AND FIN_NOTGate_0 = FIN_ANDGate_156 AND FIN_NOTGate_0 = FIN_ANDGate_157 AND FIN_NOTGate_0 = FIN_ANDGate_158 AND FIN_NOTGate_0 = FIN_ANDGate_159 AND FIN_NOTGate_0 = FIN_ANDGate_160 AND FIN_NOTGate_0 = FIN_ANDGate_161 AND FIN_NOTGate_0 = FIN_ANDGate_162 AND FIN_NOTGate_0 = FIN_ANDGate_163 AND FIN_NOTGate_0 = FIN_ANDGate_164 AND FIN_NOTGate_0 = FIN_ANDGate_165 AND FIN_NOTGate_0 = FIN_ANDGate_166 AND FIN_NOTGate_0 = FIN_ANDGate_167 AND FIN_NOTGate_0 = FIN_ANDGate_168 AND FIN_NOTGate_0 = FIN_ANDGate_169 AND FIN_NOTGate_0 = FIN_ANDGate_170 AND FIN_NOTGate_0 = FIN_ANDGate_171 AND FIN_NOTGate_0 = FIN_ANDGate_172 AND FIN_NOTGate_0 = FIN_ANDGate_173 AND FIN_NOTGate_0 = FIN_ANDGate_174 AND FIN_NOTGate_0 = FIN_ANDGate_175 AND FIN_NOTGate_0 = FIN_ANDGate_176 AND FIN_NOTGate_0 = FIN_ANDGate_177 AND FIN_NOTGate_0 = FIN_ANDGate_178 AND FIN_NOTGate_0 = FIN_ANDGate_179 AND FIN_NOTGate_0 = FIN_ANDGate_180 AND FIN_NOTGate_0 = FIN_ANDGate_181 AND FIN_NOTGate_0 = FIN_ANDGate_182 AND FIN_NOTGate_0 = FIN_ANDGate_183 AND FIN_NOTGate_0 = FIN_ANDGate_184 AND FIN_NOTGate_0 = FIN_ANDGate_185 AND FIN_NOTGate_0 = FIN_ANDGate_186 AND FIN_NOTGate_0 = FIN_ANDGate_187 AND FIN_NOTGate_0 = FIN_ANDGate_188 AND FIN_NOTGate_0 = FIN_ANDGate_189 AND FIN_NOTGate_0 = FIN_ANDGate_190 AND FIN_NOTGate_0 = FIN_ANDGate_191 AND FIN_NOTGate_0 = FIN_ANDGate_192 AND FIN_NOTGate_0 = FIN_ANDGate_193 AND FIN_NOTGate_0 = FIN_ANDGate_194 AND FIN_NOTGate_0 = FIN_ANDGate_195 AND FIN_NOTGate_0 = FIN_ANDGate_196 AND FIN_NOTGate_0 = FIN_ANDGate_197 AND FIN_NOTGate_0 = FIN_ANDGate_198 AND FIN_NOTGate_0 = FIN_ANDGate_199 AND FIN_NOTGate_0 = FIN_ANDGate_200 AND FIN_NOTGate_0 = FIN_ANDGate_201 AND FIN_NOTGate_0 = FIN_ANDGate_202 AND FIN_NOTGate_0 = FIN_ANDGate_203 AND FIN_NOTGate_0 = FIN_ANDGate_204 AND FIN_NOTGate_0 = FIN_ANDGate_205 AND FIN_NOTGate_0 = FIN_ANDGate_206 AND FIN_NOTGate_0 = FIN_ANDGate_207 AND FIN_NOTGate_0 = FIN_ANDGate_208 AND FIN_NOTGate_0 = FIN_ANDGate_209 AND FIN_NOTGate_0 = FIN_ANDGate_210 AND FIN_NOTGate_0 = FIN_ANDGate_211 AND FIN_NOTGate_0 = FIN_ANDGate_212 AND FIN_NOTGate_0 = FIN_ANDGate_213 AND FIN_NOTGate_0 = FIN_ANDGate_214 AND FIN_NOTGate_0 = FIN_ANDGate_215 AND FIN_NOTGate_0 = FIN_ANDGate_216 AND FIN_NOTGate_0 = FIN_ANDGate_217 AND FIN_NOTGate_0 = FIN_ANDGate_218 AND FIN_NOTGate_0 = FIN_ANDGate_219 AND FIN_NOTGate_0 = FIN_ANDGate_220 AND FIN_NOTGate_0 = FIN_ANDGate_221 AND FIN_NOTGate_0 = FIN_ANDGate_222 AND FIN_NOTGate_0 = FIN_ANDGate_223 AND FIN_NOTGate_0 = FIN_ANDGate_224 AND FIN_NOTGate_0 = FIN_ANDGate_225 AND FIN_NOTGate_0 = FIN_ANDGate_226 AND FIN_NOTGate_0 = FIN_ANDGate_227 AND FIN_NOTGate_0 = FIN_ANDGate_228 AND FIN_NOTGate_0 = FIN_ANDGate_229 AND FIN_NOTGate_0 = FIN_ANDGate_230 AND FIN_NOTGate_0 = FIN_ANDGate_231 AND FIN_NOTGate_0 = FIN_ANDGate_232 AND FIN_NOTGate_0 = FIN_ANDGate_233 AND FIN_NOTGate_0 = FIN_ANDGate_234 AND FIN_NOTGate_0 = FIN_ANDGate_235 AND FIN_NOTGate_0 = FIN_ANDGate_236 AND FIN_NOTGate_0 = FIN_ANDGate_237 AND FIN_NOTGate_0 = FIN_ANDGate_238 AND FIN_NOTGate_0 = FIN_ANDGate_239 AND FIN_NOTGate_0 = FIN_ANDGate_240 AND FIN_NOTGate_0 = FIN_ANDGate_241 AND FIN_NOTGate_0 = FIN_ANDGate_242 AND FIN_NOTGate_0 = FIN_ANDGate_243 AND FIN_NOTGate_0 = FIN_ANDGate_244 AND FIN_NOTGate_0 = FIN_ANDGate_245 AND FIN_NOTGate_0 = FIN_ANDGate_246 AND FIN_NOTGate_0 = FIN_ANDGate_247 AND FIN_NOTGate_0 = FIN_ANDGate_248 AND FIN_NOTGate_0 = FIN_ANDGate_249 AND FIN_NOTGate_0 = FIN_ANDGate_250 AND FIN_NOTGate_0 = FIN_ANDGate_251 AND FIN_NOTGate_0 = FIN_ANDGate_252 AND FIN_NOTGate_0 = FIN_ANDGate_253 AND FIN_NOTGate_0 = FIN_ANDGate_254 AND FIN_NOTGate_0 = FIN_ANDGate_255 then
        FIN <= FIN_NOTGate_0;
      end if;
    end process;

    -- Propagate all clocked and feedback signals
    process(
        CLK,
        RST)

        variable readyflag: std_logic;
    begin
        if RST = '1' then
            RDY <= '0';
            readyflag := '1';
        elsif rising_edge(CLK) then
            if ENB = '1' then
                readyflag := not readyflag;
                RDY <= readyflag;


            end if;
        end if;
    end process;



-- User defined processes here
-- #### USER-DATA-CODE-START
-- #### USER-DATA-CODE-END

end RTL;