library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- library SYSTEM_TYPES;
use work.SYSTEM_TYPES.ALL;

-- library CUSTOM_TYPES;
use work.CUSTOM_TYPES.ALL;

-- User defined packages here
-- #### USER-DATA-IMPORTS-START
-- #### USER-DATA-IMPORTS-END

entity Decoder_n_Bit_export is
  port(

    -- Top-level bus DecoderInput_0 signals
    DecoderInput_0_Value: in STD_LOGIC;

    -- Top-level bus DecoderNOTInput_0 signals
    DecoderNOTInput_0_Value: out STD_LOGIC;

    -- Top-level bus DecoderInput_1 signals
    DecoderInput_1_Value: in STD_LOGIC;

    -- Top-level bus DecoderNOTInput_1 signals
    DecoderNOTInput_1_Value: out STD_LOGIC;

    -- Top-level bus DecoderInput_2 signals
    DecoderInput_2_Value: in STD_LOGIC;

    -- Top-level bus DecoderNOTInput_2 signals
    DecoderNOTInput_2_Value: out STD_LOGIC;

    -- Top-level bus DecoderInput_3 signals
    DecoderInput_3_Value: in STD_LOGIC;

    -- Top-level bus DecoderNOTInput_3 signals
    DecoderNOTInput_3_Value: out STD_LOGIC;

    -- Top-level bus DecoderInput_4 signals
    DecoderInput_4_Value: in STD_LOGIC;

    -- Top-level bus DecoderNOTInput_4 signals
    DecoderNOTInput_4_Value: out STD_LOGIC;

    -- Top-level bus DecoderInput_5 signals
    DecoderInput_5_Value: in STD_LOGIC;

    -- Top-level bus DecoderNOTInput_5 signals
    DecoderNOTInput_5_Value: out STD_LOGIC;

    -- Top-level bus DecoderInput_6 signals
    DecoderInput_6_Value: in STD_LOGIC;

    -- Top-level bus DecoderNOTInput_6 signals
    DecoderNOTInput_6_Value: out STD_LOGIC;

    -- Top-level bus DecoderInput_7 signals
    DecoderInput_7_Value: in STD_LOGIC;

    -- Top-level bus DecoderNOTInput_7 signals
    DecoderNOTInput_7_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_0 signals
    DecoderOutput_0_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_1 signals
    DecoderOutput_1_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_2 signals
    DecoderOutput_2_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_3 signals
    DecoderOutput_3_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_4 signals
    DecoderOutput_4_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_5 signals
    DecoderOutput_5_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_6 signals
    DecoderOutput_6_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_7 signals
    DecoderOutput_7_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_8 signals
    DecoderOutput_8_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_9 signals
    DecoderOutput_9_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_10 signals
    DecoderOutput_10_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_11 signals
    DecoderOutput_11_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_12 signals
    DecoderOutput_12_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_13 signals
    DecoderOutput_13_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_14 signals
    DecoderOutput_14_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_15 signals
    DecoderOutput_15_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_16 signals
    DecoderOutput_16_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_17 signals
    DecoderOutput_17_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_18 signals
    DecoderOutput_18_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_19 signals
    DecoderOutput_19_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_20 signals
    DecoderOutput_20_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_21 signals
    DecoderOutput_21_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_22 signals
    DecoderOutput_22_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_23 signals
    DecoderOutput_23_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_24 signals
    DecoderOutput_24_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_25 signals
    DecoderOutput_25_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_26 signals
    DecoderOutput_26_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_27 signals
    DecoderOutput_27_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_28 signals
    DecoderOutput_28_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_29 signals
    DecoderOutput_29_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_30 signals
    DecoderOutput_30_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_31 signals
    DecoderOutput_31_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_32 signals
    DecoderOutput_32_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_33 signals
    DecoderOutput_33_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_34 signals
    DecoderOutput_34_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_35 signals
    DecoderOutput_35_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_36 signals
    DecoderOutput_36_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_37 signals
    DecoderOutput_37_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_38 signals
    DecoderOutput_38_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_39 signals
    DecoderOutput_39_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_40 signals
    DecoderOutput_40_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_41 signals
    DecoderOutput_41_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_42 signals
    DecoderOutput_42_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_43 signals
    DecoderOutput_43_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_44 signals
    DecoderOutput_44_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_45 signals
    DecoderOutput_45_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_46 signals
    DecoderOutput_46_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_47 signals
    DecoderOutput_47_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_48 signals
    DecoderOutput_48_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_49 signals
    DecoderOutput_49_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_50 signals
    DecoderOutput_50_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_51 signals
    DecoderOutput_51_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_52 signals
    DecoderOutput_52_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_53 signals
    DecoderOutput_53_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_54 signals
    DecoderOutput_54_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_55 signals
    DecoderOutput_55_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_56 signals
    DecoderOutput_56_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_57 signals
    DecoderOutput_57_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_58 signals
    DecoderOutput_58_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_59 signals
    DecoderOutput_59_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_60 signals
    DecoderOutput_60_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_61 signals
    DecoderOutput_61_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_62 signals
    DecoderOutput_62_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_63 signals
    DecoderOutput_63_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_64 signals
    DecoderOutput_64_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_65 signals
    DecoderOutput_65_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_66 signals
    DecoderOutput_66_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_67 signals
    DecoderOutput_67_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_68 signals
    DecoderOutput_68_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_69 signals
    DecoderOutput_69_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_70 signals
    DecoderOutput_70_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_71 signals
    DecoderOutput_71_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_72 signals
    DecoderOutput_72_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_73 signals
    DecoderOutput_73_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_74 signals
    DecoderOutput_74_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_75 signals
    DecoderOutput_75_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_76 signals
    DecoderOutput_76_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_77 signals
    DecoderOutput_77_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_78 signals
    DecoderOutput_78_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_79 signals
    DecoderOutput_79_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_80 signals
    DecoderOutput_80_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_81 signals
    DecoderOutput_81_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_82 signals
    DecoderOutput_82_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_83 signals
    DecoderOutput_83_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_84 signals
    DecoderOutput_84_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_85 signals
    DecoderOutput_85_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_86 signals
    DecoderOutput_86_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_87 signals
    DecoderOutput_87_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_88 signals
    DecoderOutput_88_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_89 signals
    DecoderOutput_89_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_90 signals
    DecoderOutput_90_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_91 signals
    DecoderOutput_91_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_92 signals
    DecoderOutput_92_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_93 signals
    DecoderOutput_93_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_94 signals
    DecoderOutput_94_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_95 signals
    DecoderOutput_95_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_96 signals
    DecoderOutput_96_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_97 signals
    DecoderOutput_97_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_98 signals
    DecoderOutput_98_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_99 signals
    DecoderOutput_99_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_100 signals
    DecoderOutput_100_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_101 signals
    DecoderOutput_101_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_102 signals
    DecoderOutput_102_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_103 signals
    DecoderOutput_103_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_104 signals
    DecoderOutput_104_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_105 signals
    DecoderOutput_105_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_106 signals
    DecoderOutput_106_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_107 signals
    DecoderOutput_107_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_108 signals
    DecoderOutput_108_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_109 signals
    DecoderOutput_109_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_110 signals
    DecoderOutput_110_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_111 signals
    DecoderOutput_111_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_112 signals
    DecoderOutput_112_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_113 signals
    DecoderOutput_113_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_114 signals
    DecoderOutput_114_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_115 signals
    DecoderOutput_115_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_116 signals
    DecoderOutput_116_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_117 signals
    DecoderOutput_117_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_118 signals
    DecoderOutput_118_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_119 signals
    DecoderOutput_119_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_120 signals
    DecoderOutput_120_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_121 signals
    DecoderOutput_121_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_122 signals
    DecoderOutput_122_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_123 signals
    DecoderOutput_123_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_124 signals
    DecoderOutput_124_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_125 signals
    DecoderOutput_125_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_126 signals
    DecoderOutput_126_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_127 signals
    DecoderOutput_127_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_128 signals
    DecoderOutput_128_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_129 signals
    DecoderOutput_129_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_130 signals
    DecoderOutput_130_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_131 signals
    DecoderOutput_131_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_132 signals
    DecoderOutput_132_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_133 signals
    DecoderOutput_133_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_134 signals
    DecoderOutput_134_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_135 signals
    DecoderOutput_135_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_136 signals
    DecoderOutput_136_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_137 signals
    DecoderOutput_137_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_138 signals
    DecoderOutput_138_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_139 signals
    DecoderOutput_139_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_140 signals
    DecoderOutput_140_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_141 signals
    DecoderOutput_141_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_142 signals
    DecoderOutput_142_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_143 signals
    DecoderOutput_143_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_144 signals
    DecoderOutput_144_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_145 signals
    DecoderOutput_145_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_146 signals
    DecoderOutput_146_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_147 signals
    DecoderOutput_147_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_148 signals
    DecoderOutput_148_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_149 signals
    DecoderOutput_149_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_150 signals
    DecoderOutput_150_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_151 signals
    DecoderOutput_151_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_152 signals
    DecoderOutput_152_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_153 signals
    DecoderOutput_153_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_154 signals
    DecoderOutput_154_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_155 signals
    DecoderOutput_155_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_156 signals
    DecoderOutput_156_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_157 signals
    DecoderOutput_157_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_158 signals
    DecoderOutput_158_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_159 signals
    DecoderOutput_159_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_160 signals
    DecoderOutput_160_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_161 signals
    DecoderOutput_161_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_162 signals
    DecoderOutput_162_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_163 signals
    DecoderOutput_163_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_164 signals
    DecoderOutput_164_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_165 signals
    DecoderOutput_165_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_166 signals
    DecoderOutput_166_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_167 signals
    DecoderOutput_167_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_168 signals
    DecoderOutput_168_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_169 signals
    DecoderOutput_169_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_170 signals
    DecoderOutput_170_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_171 signals
    DecoderOutput_171_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_172 signals
    DecoderOutput_172_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_173 signals
    DecoderOutput_173_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_174 signals
    DecoderOutput_174_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_175 signals
    DecoderOutput_175_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_176 signals
    DecoderOutput_176_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_177 signals
    DecoderOutput_177_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_178 signals
    DecoderOutput_178_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_179 signals
    DecoderOutput_179_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_180 signals
    DecoderOutput_180_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_181 signals
    DecoderOutput_181_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_182 signals
    DecoderOutput_182_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_183 signals
    DecoderOutput_183_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_184 signals
    DecoderOutput_184_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_185 signals
    DecoderOutput_185_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_186 signals
    DecoderOutput_186_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_187 signals
    DecoderOutput_187_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_188 signals
    DecoderOutput_188_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_189 signals
    DecoderOutput_189_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_190 signals
    DecoderOutput_190_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_191 signals
    DecoderOutput_191_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_192 signals
    DecoderOutput_192_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_193 signals
    DecoderOutput_193_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_194 signals
    DecoderOutput_194_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_195 signals
    DecoderOutput_195_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_196 signals
    DecoderOutput_196_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_197 signals
    DecoderOutput_197_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_198 signals
    DecoderOutput_198_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_199 signals
    DecoderOutput_199_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_200 signals
    DecoderOutput_200_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_201 signals
    DecoderOutput_201_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_202 signals
    DecoderOutput_202_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_203 signals
    DecoderOutput_203_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_204 signals
    DecoderOutput_204_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_205 signals
    DecoderOutput_205_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_206 signals
    DecoderOutput_206_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_207 signals
    DecoderOutput_207_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_208 signals
    DecoderOutput_208_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_209 signals
    DecoderOutput_209_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_210 signals
    DecoderOutput_210_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_211 signals
    DecoderOutput_211_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_212 signals
    DecoderOutput_212_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_213 signals
    DecoderOutput_213_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_214 signals
    DecoderOutput_214_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_215 signals
    DecoderOutput_215_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_216 signals
    DecoderOutput_216_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_217 signals
    DecoderOutput_217_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_218 signals
    DecoderOutput_218_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_219 signals
    DecoderOutput_219_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_220 signals
    DecoderOutput_220_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_221 signals
    DecoderOutput_221_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_222 signals
    DecoderOutput_222_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_223 signals
    DecoderOutput_223_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_224 signals
    DecoderOutput_224_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_225 signals
    DecoderOutput_225_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_226 signals
    DecoderOutput_226_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_227 signals
    DecoderOutput_227_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_228 signals
    DecoderOutput_228_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_229 signals
    DecoderOutput_229_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_230 signals
    DecoderOutput_230_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_231 signals
    DecoderOutput_231_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_232 signals
    DecoderOutput_232_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_233 signals
    DecoderOutput_233_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_234 signals
    DecoderOutput_234_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_235 signals
    DecoderOutput_235_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_236 signals
    DecoderOutput_236_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_237 signals
    DecoderOutput_237_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_238 signals
    DecoderOutput_238_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_239 signals
    DecoderOutput_239_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_240 signals
    DecoderOutput_240_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_241 signals
    DecoderOutput_241_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_242 signals
    DecoderOutput_242_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_243 signals
    DecoderOutput_243_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_244 signals
    DecoderOutput_244_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_245 signals
    DecoderOutput_245_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_246 signals
    DecoderOutput_246_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_247 signals
    DecoderOutput_247_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_248 signals
    DecoderOutput_248_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_249 signals
    DecoderOutput_249_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_250 signals
    DecoderOutput_250_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_251 signals
    DecoderOutput_251_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_252 signals
    DecoderOutput_252_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_253 signals
    DecoderOutput_253_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_254 signals
    DecoderOutput_254_Value: out STD_LOGIC;

    -- Top-level bus DecoderOutput_255 signals
    DecoderOutput_255_Value: out STD_LOGIC;


    -- User defined signals here
    -- #### USER-DATA-ENTITYSIGNALS-START
    -- #### USER-DATA-ENTITYSIGNALS-END


    -- Enable signal
    ENB : in STD_LOGIC;

	-- Reset signal
    RST : in STD_LOGIC;

    -- Finished signal
    FIN : out Std_logic;

    -- Clock signal
    CLK : in STD_LOGIC
  );
end Decoder_n_Bit_export;



architecture RTL of Decoder_n_Bit_export is  
  -- User defined signals here
  -- #### USER-DATA-SIGNALS-START
  -- #### USER-DATA-SIGNALS-END


begin

    -- Entity Decoder_n_Bit signals
    Decoder_n_Bit: entity work.Decoder_n_Bit
    port map (
        -- Input bus DecoderInput_0
        DecoderInput_0_Value => DecoderInput_0_Value,

        -- Output bus DecoderNOTInput_0
        DecoderNOTInput_0_Value => DecoderNOTInput_0_Value,

        -- Input bus DecoderInput_1
        DecoderInput_1_Value => DecoderInput_1_Value,

        -- Output bus DecoderNOTInput_1
        DecoderNOTInput_1_Value => DecoderNOTInput_1_Value,

        -- Input bus DecoderInput_2
        DecoderInput_2_Value => DecoderInput_2_Value,

        -- Output bus DecoderNOTInput_2
        DecoderNOTInput_2_Value => DecoderNOTInput_2_Value,

        -- Input bus DecoderInput_3
        DecoderInput_3_Value => DecoderInput_3_Value,

        -- Output bus DecoderNOTInput_3
        DecoderNOTInput_3_Value => DecoderNOTInput_3_Value,

        -- Input bus DecoderInput_4
        DecoderInput_4_Value => DecoderInput_4_Value,

        -- Output bus DecoderNOTInput_4
        DecoderNOTInput_4_Value => DecoderNOTInput_4_Value,

        -- Input bus DecoderInput_5
        DecoderInput_5_Value => DecoderInput_5_Value,

        -- Output bus DecoderNOTInput_5
        DecoderNOTInput_5_Value => DecoderNOTInput_5_Value,

        -- Input bus DecoderInput_6
        DecoderInput_6_Value => DecoderInput_6_Value,

        -- Output bus DecoderNOTInput_6
        DecoderNOTInput_6_Value => DecoderNOTInput_6_Value,

        -- Input bus DecoderInput_7
        DecoderInput_7_Value => DecoderInput_7_Value,

        -- Output bus DecoderNOTInput_7
        DecoderNOTInput_7_Value => DecoderNOTInput_7_Value,

        -- Output bus DecoderOutput_0
        DecoderOutput_0_Value => DecoderOutput_0_Value,

        -- Output bus DecoderOutput_1
        DecoderOutput_1_Value => DecoderOutput_1_Value,

        -- Output bus DecoderOutput_2
        DecoderOutput_2_Value => DecoderOutput_2_Value,

        -- Output bus DecoderOutput_3
        DecoderOutput_3_Value => DecoderOutput_3_Value,

        -- Output bus DecoderOutput_4
        DecoderOutput_4_Value => DecoderOutput_4_Value,

        -- Output bus DecoderOutput_5
        DecoderOutput_5_Value => DecoderOutput_5_Value,

        -- Output bus DecoderOutput_6
        DecoderOutput_6_Value => DecoderOutput_6_Value,

        -- Output bus DecoderOutput_7
        DecoderOutput_7_Value => DecoderOutput_7_Value,

        -- Output bus DecoderOutput_8
        DecoderOutput_8_Value => DecoderOutput_8_Value,

        -- Output bus DecoderOutput_9
        DecoderOutput_9_Value => DecoderOutput_9_Value,

        -- Output bus DecoderOutput_10
        DecoderOutput_10_Value => DecoderOutput_10_Value,

        -- Output bus DecoderOutput_11
        DecoderOutput_11_Value => DecoderOutput_11_Value,

        -- Output bus DecoderOutput_12
        DecoderOutput_12_Value => DecoderOutput_12_Value,

        -- Output bus DecoderOutput_13
        DecoderOutput_13_Value => DecoderOutput_13_Value,

        -- Output bus DecoderOutput_14
        DecoderOutput_14_Value => DecoderOutput_14_Value,

        -- Output bus DecoderOutput_15
        DecoderOutput_15_Value => DecoderOutput_15_Value,

        -- Output bus DecoderOutput_16
        DecoderOutput_16_Value => DecoderOutput_16_Value,

        -- Output bus DecoderOutput_17
        DecoderOutput_17_Value => DecoderOutput_17_Value,

        -- Output bus DecoderOutput_18
        DecoderOutput_18_Value => DecoderOutput_18_Value,

        -- Output bus DecoderOutput_19
        DecoderOutput_19_Value => DecoderOutput_19_Value,

        -- Output bus DecoderOutput_20
        DecoderOutput_20_Value => DecoderOutput_20_Value,

        -- Output bus DecoderOutput_21
        DecoderOutput_21_Value => DecoderOutput_21_Value,

        -- Output bus DecoderOutput_22
        DecoderOutput_22_Value => DecoderOutput_22_Value,

        -- Output bus DecoderOutput_23
        DecoderOutput_23_Value => DecoderOutput_23_Value,

        -- Output bus DecoderOutput_24
        DecoderOutput_24_Value => DecoderOutput_24_Value,

        -- Output bus DecoderOutput_25
        DecoderOutput_25_Value => DecoderOutput_25_Value,

        -- Output bus DecoderOutput_26
        DecoderOutput_26_Value => DecoderOutput_26_Value,

        -- Output bus DecoderOutput_27
        DecoderOutput_27_Value => DecoderOutput_27_Value,

        -- Output bus DecoderOutput_28
        DecoderOutput_28_Value => DecoderOutput_28_Value,

        -- Output bus DecoderOutput_29
        DecoderOutput_29_Value => DecoderOutput_29_Value,

        -- Output bus DecoderOutput_30
        DecoderOutput_30_Value => DecoderOutput_30_Value,

        -- Output bus DecoderOutput_31
        DecoderOutput_31_Value => DecoderOutput_31_Value,

        -- Output bus DecoderOutput_32
        DecoderOutput_32_Value => DecoderOutput_32_Value,

        -- Output bus DecoderOutput_33
        DecoderOutput_33_Value => DecoderOutput_33_Value,

        -- Output bus DecoderOutput_34
        DecoderOutput_34_Value => DecoderOutput_34_Value,

        -- Output bus DecoderOutput_35
        DecoderOutput_35_Value => DecoderOutput_35_Value,

        -- Output bus DecoderOutput_36
        DecoderOutput_36_Value => DecoderOutput_36_Value,

        -- Output bus DecoderOutput_37
        DecoderOutput_37_Value => DecoderOutput_37_Value,

        -- Output bus DecoderOutput_38
        DecoderOutput_38_Value => DecoderOutput_38_Value,

        -- Output bus DecoderOutput_39
        DecoderOutput_39_Value => DecoderOutput_39_Value,

        -- Output bus DecoderOutput_40
        DecoderOutput_40_Value => DecoderOutput_40_Value,

        -- Output bus DecoderOutput_41
        DecoderOutput_41_Value => DecoderOutput_41_Value,

        -- Output bus DecoderOutput_42
        DecoderOutput_42_Value => DecoderOutput_42_Value,

        -- Output bus DecoderOutput_43
        DecoderOutput_43_Value => DecoderOutput_43_Value,

        -- Output bus DecoderOutput_44
        DecoderOutput_44_Value => DecoderOutput_44_Value,

        -- Output bus DecoderOutput_45
        DecoderOutput_45_Value => DecoderOutput_45_Value,

        -- Output bus DecoderOutput_46
        DecoderOutput_46_Value => DecoderOutput_46_Value,

        -- Output bus DecoderOutput_47
        DecoderOutput_47_Value => DecoderOutput_47_Value,

        -- Output bus DecoderOutput_48
        DecoderOutput_48_Value => DecoderOutput_48_Value,

        -- Output bus DecoderOutput_49
        DecoderOutput_49_Value => DecoderOutput_49_Value,

        -- Output bus DecoderOutput_50
        DecoderOutput_50_Value => DecoderOutput_50_Value,

        -- Output bus DecoderOutput_51
        DecoderOutput_51_Value => DecoderOutput_51_Value,

        -- Output bus DecoderOutput_52
        DecoderOutput_52_Value => DecoderOutput_52_Value,

        -- Output bus DecoderOutput_53
        DecoderOutput_53_Value => DecoderOutput_53_Value,

        -- Output bus DecoderOutput_54
        DecoderOutput_54_Value => DecoderOutput_54_Value,

        -- Output bus DecoderOutput_55
        DecoderOutput_55_Value => DecoderOutput_55_Value,

        -- Output bus DecoderOutput_56
        DecoderOutput_56_Value => DecoderOutput_56_Value,

        -- Output bus DecoderOutput_57
        DecoderOutput_57_Value => DecoderOutput_57_Value,

        -- Output bus DecoderOutput_58
        DecoderOutput_58_Value => DecoderOutput_58_Value,

        -- Output bus DecoderOutput_59
        DecoderOutput_59_Value => DecoderOutput_59_Value,

        -- Output bus DecoderOutput_60
        DecoderOutput_60_Value => DecoderOutput_60_Value,

        -- Output bus DecoderOutput_61
        DecoderOutput_61_Value => DecoderOutput_61_Value,

        -- Output bus DecoderOutput_62
        DecoderOutput_62_Value => DecoderOutput_62_Value,

        -- Output bus DecoderOutput_63
        DecoderOutput_63_Value => DecoderOutput_63_Value,

        -- Output bus DecoderOutput_64
        DecoderOutput_64_Value => DecoderOutput_64_Value,

        -- Output bus DecoderOutput_65
        DecoderOutput_65_Value => DecoderOutput_65_Value,

        -- Output bus DecoderOutput_66
        DecoderOutput_66_Value => DecoderOutput_66_Value,

        -- Output bus DecoderOutput_67
        DecoderOutput_67_Value => DecoderOutput_67_Value,

        -- Output bus DecoderOutput_68
        DecoderOutput_68_Value => DecoderOutput_68_Value,

        -- Output bus DecoderOutput_69
        DecoderOutput_69_Value => DecoderOutput_69_Value,

        -- Output bus DecoderOutput_70
        DecoderOutput_70_Value => DecoderOutput_70_Value,

        -- Output bus DecoderOutput_71
        DecoderOutput_71_Value => DecoderOutput_71_Value,

        -- Output bus DecoderOutput_72
        DecoderOutput_72_Value => DecoderOutput_72_Value,

        -- Output bus DecoderOutput_73
        DecoderOutput_73_Value => DecoderOutput_73_Value,

        -- Output bus DecoderOutput_74
        DecoderOutput_74_Value => DecoderOutput_74_Value,

        -- Output bus DecoderOutput_75
        DecoderOutput_75_Value => DecoderOutput_75_Value,

        -- Output bus DecoderOutput_76
        DecoderOutput_76_Value => DecoderOutput_76_Value,

        -- Output bus DecoderOutput_77
        DecoderOutput_77_Value => DecoderOutput_77_Value,

        -- Output bus DecoderOutput_78
        DecoderOutput_78_Value => DecoderOutput_78_Value,

        -- Output bus DecoderOutput_79
        DecoderOutput_79_Value => DecoderOutput_79_Value,

        -- Output bus DecoderOutput_80
        DecoderOutput_80_Value => DecoderOutput_80_Value,

        -- Output bus DecoderOutput_81
        DecoderOutput_81_Value => DecoderOutput_81_Value,

        -- Output bus DecoderOutput_82
        DecoderOutput_82_Value => DecoderOutput_82_Value,

        -- Output bus DecoderOutput_83
        DecoderOutput_83_Value => DecoderOutput_83_Value,

        -- Output bus DecoderOutput_84
        DecoderOutput_84_Value => DecoderOutput_84_Value,

        -- Output bus DecoderOutput_85
        DecoderOutput_85_Value => DecoderOutput_85_Value,

        -- Output bus DecoderOutput_86
        DecoderOutput_86_Value => DecoderOutput_86_Value,

        -- Output bus DecoderOutput_87
        DecoderOutput_87_Value => DecoderOutput_87_Value,

        -- Output bus DecoderOutput_88
        DecoderOutput_88_Value => DecoderOutput_88_Value,

        -- Output bus DecoderOutput_89
        DecoderOutput_89_Value => DecoderOutput_89_Value,

        -- Output bus DecoderOutput_90
        DecoderOutput_90_Value => DecoderOutput_90_Value,

        -- Output bus DecoderOutput_91
        DecoderOutput_91_Value => DecoderOutput_91_Value,

        -- Output bus DecoderOutput_92
        DecoderOutput_92_Value => DecoderOutput_92_Value,

        -- Output bus DecoderOutput_93
        DecoderOutput_93_Value => DecoderOutput_93_Value,

        -- Output bus DecoderOutput_94
        DecoderOutput_94_Value => DecoderOutput_94_Value,

        -- Output bus DecoderOutput_95
        DecoderOutput_95_Value => DecoderOutput_95_Value,

        -- Output bus DecoderOutput_96
        DecoderOutput_96_Value => DecoderOutput_96_Value,

        -- Output bus DecoderOutput_97
        DecoderOutput_97_Value => DecoderOutput_97_Value,

        -- Output bus DecoderOutput_98
        DecoderOutput_98_Value => DecoderOutput_98_Value,

        -- Output bus DecoderOutput_99
        DecoderOutput_99_Value => DecoderOutput_99_Value,

        -- Output bus DecoderOutput_100
        DecoderOutput_100_Value => DecoderOutput_100_Value,

        -- Output bus DecoderOutput_101
        DecoderOutput_101_Value => DecoderOutput_101_Value,

        -- Output bus DecoderOutput_102
        DecoderOutput_102_Value => DecoderOutput_102_Value,

        -- Output bus DecoderOutput_103
        DecoderOutput_103_Value => DecoderOutput_103_Value,

        -- Output bus DecoderOutput_104
        DecoderOutput_104_Value => DecoderOutput_104_Value,

        -- Output bus DecoderOutput_105
        DecoderOutput_105_Value => DecoderOutput_105_Value,

        -- Output bus DecoderOutput_106
        DecoderOutput_106_Value => DecoderOutput_106_Value,

        -- Output bus DecoderOutput_107
        DecoderOutput_107_Value => DecoderOutput_107_Value,

        -- Output bus DecoderOutput_108
        DecoderOutput_108_Value => DecoderOutput_108_Value,

        -- Output bus DecoderOutput_109
        DecoderOutput_109_Value => DecoderOutput_109_Value,

        -- Output bus DecoderOutput_110
        DecoderOutput_110_Value => DecoderOutput_110_Value,

        -- Output bus DecoderOutput_111
        DecoderOutput_111_Value => DecoderOutput_111_Value,

        -- Output bus DecoderOutput_112
        DecoderOutput_112_Value => DecoderOutput_112_Value,

        -- Output bus DecoderOutput_113
        DecoderOutput_113_Value => DecoderOutput_113_Value,

        -- Output bus DecoderOutput_114
        DecoderOutput_114_Value => DecoderOutput_114_Value,

        -- Output bus DecoderOutput_115
        DecoderOutput_115_Value => DecoderOutput_115_Value,

        -- Output bus DecoderOutput_116
        DecoderOutput_116_Value => DecoderOutput_116_Value,

        -- Output bus DecoderOutput_117
        DecoderOutput_117_Value => DecoderOutput_117_Value,

        -- Output bus DecoderOutput_118
        DecoderOutput_118_Value => DecoderOutput_118_Value,

        -- Output bus DecoderOutput_119
        DecoderOutput_119_Value => DecoderOutput_119_Value,

        -- Output bus DecoderOutput_120
        DecoderOutput_120_Value => DecoderOutput_120_Value,

        -- Output bus DecoderOutput_121
        DecoderOutput_121_Value => DecoderOutput_121_Value,

        -- Output bus DecoderOutput_122
        DecoderOutput_122_Value => DecoderOutput_122_Value,

        -- Output bus DecoderOutput_123
        DecoderOutput_123_Value => DecoderOutput_123_Value,

        -- Output bus DecoderOutput_124
        DecoderOutput_124_Value => DecoderOutput_124_Value,

        -- Output bus DecoderOutput_125
        DecoderOutput_125_Value => DecoderOutput_125_Value,

        -- Output bus DecoderOutput_126
        DecoderOutput_126_Value => DecoderOutput_126_Value,

        -- Output bus DecoderOutput_127
        DecoderOutput_127_Value => DecoderOutput_127_Value,

        -- Output bus DecoderOutput_128
        DecoderOutput_128_Value => DecoderOutput_128_Value,

        -- Output bus DecoderOutput_129
        DecoderOutput_129_Value => DecoderOutput_129_Value,

        -- Output bus DecoderOutput_130
        DecoderOutput_130_Value => DecoderOutput_130_Value,

        -- Output bus DecoderOutput_131
        DecoderOutput_131_Value => DecoderOutput_131_Value,

        -- Output bus DecoderOutput_132
        DecoderOutput_132_Value => DecoderOutput_132_Value,

        -- Output bus DecoderOutput_133
        DecoderOutput_133_Value => DecoderOutput_133_Value,

        -- Output bus DecoderOutput_134
        DecoderOutput_134_Value => DecoderOutput_134_Value,

        -- Output bus DecoderOutput_135
        DecoderOutput_135_Value => DecoderOutput_135_Value,

        -- Output bus DecoderOutput_136
        DecoderOutput_136_Value => DecoderOutput_136_Value,

        -- Output bus DecoderOutput_137
        DecoderOutput_137_Value => DecoderOutput_137_Value,

        -- Output bus DecoderOutput_138
        DecoderOutput_138_Value => DecoderOutput_138_Value,

        -- Output bus DecoderOutput_139
        DecoderOutput_139_Value => DecoderOutput_139_Value,

        -- Output bus DecoderOutput_140
        DecoderOutput_140_Value => DecoderOutput_140_Value,

        -- Output bus DecoderOutput_141
        DecoderOutput_141_Value => DecoderOutput_141_Value,

        -- Output bus DecoderOutput_142
        DecoderOutput_142_Value => DecoderOutput_142_Value,

        -- Output bus DecoderOutput_143
        DecoderOutput_143_Value => DecoderOutput_143_Value,

        -- Output bus DecoderOutput_144
        DecoderOutput_144_Value => DecoderOutput_144_Value,

        -- Output bus DecoderOutput_145
        DecoderOutput_145_Value => DecoderOutput_145_Value,

        -- Output bus DecoderOutput_146
        DecoderOutput_146_Value => DecoderOutput_146_Value,

        -- Output bus DecoderOutput_147
        DecoderOutput_147_Value => DecoderOutput_147_Value,

        -- Output bus DecoderOutput_148
        DecoderOutput_148_Value => DecoderOutput_148_Value,

        -- Output bus DecoderOutput_149
        DecoderOutput_149_Value => DecoderOutput_149_Value,

        -- Output bus DecoderOutput_150
        DecoderOutput_150_Value => DecoderOutput_150_Value,

        -- Output bus DecoderOutput_151
        DecoderOutput_151_Value => DecoderOutput_151_Value,

        -- Output bus DecoderOutput_152
        DecoderOutput_152_Value => DecoderOutput_152_Value,

        -- Output bus DecoderOutput_153
        DecoderOutput_153_Value => DecoderOutput_153_Value,

        -- Output bus DecoderOutput_154
        DecoderOutput_154_Value => DecoderOutput_154_Value,

        -- Output bus DecoderOutput_155
        DecoderOutput_155_Value => DecoderOutput_155_Value,

        -- Output bus DecoderOutput_156
        DecoderOutput_156_Value => DecoderOutput_156_Value,

        -- Output bus DecoderOutput_157
        DecoderOutput_157_Value => DecoderOutput_157_Value,

        -- Output bus DecoderOutput_158
        DecoderOutput_158_Value => DecoderOutput_158_Value,

        -- Output bus DecoderOutput_159
        DecoderOutput_159_Value => DecoderOutput_159_Value,

        -- Output bus DecoderOutput_160
        DecoderOutput_160_Value => DecoderOutput_160_Value,

        -- Output bus DecoderOutput_161
        DecoderOutput_161_Value => DecoderOutput_161_Value,

        -- Output bus DecoderOutput_162
        DecoderOutput_162_Value => DecoderOutput_162_Value,

        -- Output bus DecoderOutput_163
        DecoderOutput_163_Value => DecoderOutput_163_Value,

        -- Output bus DecoderOutput_164
        DecoderOutput_164_Value => DecoderOutput_164_Value,

        -- Output bus DecoderOutput_165
        DecoderOutput_165_Value => DecoderOutput_165_Value,

        -- Output bus DecoderOutput_166
        DecoderOutput_166_Value => DecoderOutput_166_Value,

        -- Output bus DecoderOutput_167
        DecoderOutput_167_Value => DecoderOutput_167_Value,

        -- Output bus DecoderOutput_168
        DecoderOutput_168_Value => DecoderOutput_168_Value,

        -- Output bus DecoderOutput_169
        DecoderOutput_169_Value => DecoderOutput_169_Value,

        -- Output bus DecoderOutput_170
        DecoderOutput_170_Value => DecoderOutput_170_Value,

        -- Output bus DecoderOutput_171
        DecoderOutput_171_Value => DecoderOutput_171_Value,

        -- Output bus DecoderOutput_172
        DecoderOutput_172_Value => DecoderOutput_172_Value,

        -- Output bus DecoderOutput_173
        DecoderOutput_173_Value => DecoderOutput_173_Value,

        -- Output bus DecoderOutput_174
        DecoderOutput_174_Value => DecoderOutput_174_Value,

        -- Output bus DecoderOutput_175
        DecoderOutput_175_Value => DecoderOutput_175_Value,

        -- Output bus DecoderOutput_176
        DecoderOutput_176_Value => DecoderOutput_176_Value,

        -- Output bus DecoderOutput_177
        DecoderOutput_177_Value => DecoderOutput_177_Value,

        -- Output bus DecoderOutput_178
        DecoderOutput_178_Value => DecoderOutput_178_Value,

        -- Output bus DecoderOutput_179
        DecoderOutput_179_Value => DecoderOutput_179_Value,

        -- Output bus DecoderOutput_180
        DecoderOutput_180_Value => DecoderOutput_180_Value,

        -- Output bus DecoderOutput_181
        DecoderOutput_181_Value => DecoderOutput_181_Value,

        -- Output bus DecoderOutput_182
        DecoderOutput_182_Value => DecoderOutput_182_Value,

        -- Output bus DecoderOutput_183
        DecoderOutput_183_Value => DecoderOutput_183_Value,

        -- Output bus DecoderOutput_184
        DecoderOutput_184_Value => DecoderOutput_184_Value,

        -- Output bus DecoderOutput_185
        DecoderOutput_185_Value => DecoderOutput_185_Value,

        -- Output bus DecoderOutput_186
        DecoderOutput_186_Value => DecoderOutput_186_Value,

        -- Output bus DecoderOutput_187
        DecoderOutput_187_Value => DecoderOutput_187_Value,

        -- Output bus DecoderOutput_188
        DecoderOutput_188_Value => DecoderOutput_188_Value,

        -- Output bus DecoderOutput_189
        DecoderOutput_189_Value => DecoderOutput_189_Value,

        -- Output bus DecoderOutput_190
        DecoderOutput_190_Value => DecoderOutput_190_Value,

        -- Output bus DecoderOutput_191
        DecoderOutput_191_Value => DecoderOutput_191_Value,

        -- Output bus DecoderOutput_192
        DecoderOutput_192_Value => DecoderOutput_192_Value,

        -- Output bus DecoderOutput_193
        DecoderOutput_193_Value => DecoderOutput_193_Value,

        -- Output bus DecoderOutput_194
        DecoderOutput_194_Value => DecoderOutput_194_Value,

        -- Output bus DecoderOutput_195
        DecoderOutput_195_Value => DecoderOutput_195_Value,

        -- Output bus DecoderOutput_196
        DecoderOutput_196_Value => DecoderOutput_196_Value,

        -- Output bus DecoderOutput_197
        DecoderOutput_197_Value => DecoderOutput_197_Value,

        -- Output bus DecoderOutput_198
        DecoderOutput_198_Value => DecoderOutput_198_Value,

        -- Output bus DecoderOutput_199
        DecoderOutput_199_Value => DecoderOutput_199_Value,

        -- Output bus DecoderOutput_200
        DecoderOutput_200_Value => DecoderOutput_200_Value,

        -- Output bus DecoderOutput_201
        DecoderOutput_201_Value => DecoderOutput_201_Value,

        -- Output bus DecoderOutput_202
        DecoderOutput_202_Value => DecoderOutput_202_Value,

        -- Output bus DecoderOutput_203
        DecoderOutput_203_Value => DecoderOutput_203_Value,

        -- Output bus DecoderOutput_204
        DecoderOutput_204_Value => DecoderOutput_204_Value,

        -- Output bus DecoderOutput_205
        DecoderOutput_205_Value => DecoderOutput_205_Value,

        -- Output bus DecoderOutput_206
        DecoderOutput_206_Value => DecoderOutput_206_Value,

        -- Output bus DecoderOutput_207
        DecoderOutput_207_Value => DecoderOutput_207_Value,

        -- Output bus DecoderOutput_208
        DecoderOutput_208_Value => DecoderOutput_208_Value,

        -- Output bus DecoderOutput_209
        DecoderOutput_209_Value => DecoderOutput_209_Value,

        -- Output bus DecoderOutput_210
        DecoderOutput_210_Value => DecoderOutput_210_Value,

        -- Output bus DecoderOutput_211
        DecoderOutput_211_Value => DecoderOutput_211_Value,

        -- Output bus DecoderOutput_212
        DecoderOutput_212_Value => DecoderOutput_212_Value,

        -- Output bus DecoderOutput_213
        DecoderOutput_213_Value => DecoderOutput_213_Value,

        -- Output bus DecoderOutput_214
        DecoderOutput_214_Value => DecoderOutput_214_Value,

        -- Output bus DecoderOutput_215
        DecoderOutput_215_Value => DecoderOutput_215_Value,

        -- Output bus DecoderOutput_216
        DecoderOutput_216_Value => DecoderOutput_216_Value,

        -- Output bus DecoderOutput_217
        DecoderOutput_217_Value => DecoderOutput_217_Value,

        -- Output bus DecoderOutput_218
        DecoderOutput_218_Value => DecoderOutput_218_Value,

        -- Output bus DecoderOutput_219
        DecoderOutput_219_Value => DecoderOutput_219_Value,

        -- Output bus DecoderOutput_220
        DecoderOutput_220_Value => DecoderOutput_220_Value,

        -- Output bus DecoderOutput_221
        DecoderOutput_221_Value => DecoderOutput_221_Value,

        -- Output bus DecoderOutput_222
        DecoderOutput_222_Value => DecoderOutput_222_Value,

        -- Output bus DecoderOutput_223
        DecoderOutput_223_Value => DecoderOutput_223_Value,

        -- Output bus DecoderOutput_224
        DecoderOutput_224_Value => DecoderOutput_224_Value,

        -- Output bus DecoderOutput_225
        DecoderOutput_225_Value => DecoderOutput_225_Value,

        -- Output bus DecoderOutput_226
        DecoderOutput_226_Value => DecoderOutput_226_Value,

        -- Output bus DecoderOutput_227
        DecoderOutput_227_Value => DecoderOutput_227_Value,

        -- Output bus DecoderOutput_228
        DecoderOutput_228_Value => DecoderOutput_228_Value,

        -- Output bus DecoderOutput_229
        DecoderOutput_229_Value => DecoderOutput_229_Value,

        -- Output bus DecoderOutput_230
        DecoderOutput_230_Value => DecoderOutput_230_Value,

        -- Output bus DecoderOutput_231
        DecoderOutput_231_Value => DecoderOutput_231_Value,

        -- Output bus DecoderOutput_232
        DecoderOutput_232_Value => DecoderOutput_232_Value,

        -- Output bus DecoderOutput_233
        DecoderOutput_233_Value => DecoderOutput_233_Value,

        -- Output bus DecoderOutput_234
        DecoderOutput_234_Value => DecoderOutput_234_Value,

        -- Output bus DecoderOutput_235
        DecoderOutput_235_Value => DecoderOutput_235_Value,

        -- Output bus DecoderOutput_236
        DecoderOutput_236_Value => DecoderOutput_236_Value,

        -- Output bus DecoderOutput_237
        DecoderOutput_237_Value => DecoderOutput_237_Value,

        -- Output bus DecoderOutput_238
        DecoderOutput_238_Value => DecoderOutput_238_Value,

        -- Output bus DecoderOutput_239
        DecoderOutput_239_Value => DecoderOutput_239_Value,

        -- Output bus DecoderOutput_240
        DecoderOutput_240_Value => DecoderOutput_240_Value,

        -- Output bus DecoderOutput_241
        DecoderOutput_241_Value => DecoderOutput_241_Value,

        -- Output bus DecoderOutput_242
        DecoderOutput_242_Value => DecoderOutput_242_Value,

        -- Output bus DecoderOutput_243
        DecoderOutput_243_Value => DecoderOutput_243_Value,

        -- Output bus DecoderOutput_244
        DecoderOutput_244_Value => DecoderOutput_244_Value,

        -- Output bus DecoderOutput_245
        DecoderOutput_245_Value => DecoderOutput_245_Value,

        -- Output bus DecoderOutput_246
        DecoderOutput_246_Value => DecoderOutput_246_Value,

        -- Output bus DecoderOutput_247
        DecoderOutput_247_Value => DecoderOutput_247_Value,

        -- Output bus DecoderOutput_248
        DecoderOutput_248_Value => DecoderOutput_248_Value,

        -- Output bus DecoderOutput_249
        DecoderOutput_249_Value => DecoderOutput_249_Value,

        -- Output bus DecoderOutput_250
        DecoderOutput_250_Value => DecoderOutput_250_Value,

        -- Output bus DecoderOutput_251
        DecoderOutput_251_Value => DecoderOutput_251_Value,

        -- Output bus DecoderOutput_252
        DecoderOutput_252_Value => DecoderOutput_252_Value,

        -- Output bus DecoderOutput_253
        DecoderOutput_253_Value => DecoderOutput_253_Value,

        -- Output bus DecoderOutput_254
        DecoderOutput_254_Value => DecoderOutput_254_Value,

        -- Output bus DecoderOutput_255
        DecoderOutput_255_Value => DecoderOutput_255_Value,

        ENB => ENB,
        RST => RST,
        FIN => FIN,
        CLK => CLK
    );

-- User defined processes here
-- #### USER-DATA-CODE-START
-- #### USER-DATA-CODE-END

end RTL;